module ALU(
  input        clock,
  input        reset,
  input  [8:0] io_opcode,
  input  [3:0] io_in_a,
  input  [3:0] io_in_b,
  output [3:0] io_out_a,
  output [3:0] io_out_b,
  input        io_validin_a,
  input        io_validin_b,
  output       io_validout_a,
  output       io_validout_b
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] snapshot_a; // @[ALU.scala 25:27]
  reg [3:0] snapshot_b; // @[ALU.scala 26:27]
  reg  snapshot_valid_a; // @[ALU.scala 28:33]
  reg  snapshot_valid_b; // @[ALU.scala 29:33]
  reg [3:0] temp_result_a; // @[ALU.scala 33:30]
  reg [3:0] temp_result_b; // @[ALU.scala 34:30]
  reg  temp_valid_a; // @[ALU.scala 37:29]
  reg  temp_valid_b; // @[ALU.scala 38:29]
  wire  opcode_0 = io_opcode[0]; // @[ALU.scala 41:34]
  wire  opcode_1 = io_opcode[1]; // @[ALU.scala 41:34]
  wire  opcode_2 = io_opcode[2]; // @[ALU.scala 41:34]
  wire  opcode_3 = io_opcode[3]; // @[ALU.scala 41:34]
  wire  opcode_4 = io_opcode[4]; // @[ALU.scala 41:34]
  wire  opcode_5 = io_opcode[5]; // @[ALU.scala 41:34]
  wire  opcode_6 = io_opcode[6]; // @[ALU.scala 41:34]
  wire  opcode_7 = io_opcode[7]; // @[ALU.scala 41:34]
  wire  opcode_8 = io_opcode[8]; // @[ALU.scala 41:34]
  wire  _T_1 = ~opcode_7; // @[ALU.scala 51:39]
  wire  _T_5 = opcode_6 & opcode_5; // @[ALU.scala 52:28]
  wire  _T_26 = ~opcode_4; // @[ALU.scala 93:20]
  wire  _T_27 = ~opcode_3; // @[ALU.scala 93:41]
  wire  _T_28 = ~opcode_4 & ~opcode_3; // @[ALU.scala 93:28]
  wire [3:0] _gate_a_T = ~io_in_a; // @[ALU.scala 94:17]
  wire  _T_31 = opcode_4 & _T_27; // @[ALU.scala 98:34]
  wire [3:0] _gate_a_T_1 = ~snapshot_a; // @[ALU.scala 99:17]
  wire  _T_34 = _T_26 & opcode_3; // @[ALU.scala 103:34]
  wire [3:0] _GEN_18 = _T_26 & opcode_3 ? _gate_a_T : _gate_a_T_1; // @[ALU.scala 103:55 ALU.scala 104:14 ALU.scala 109:14]
  wire [3:0] _GEN_22 = opcode_4 & _T_27 ? _gate_a_T_1 : _GEN_18; // @[ALU.scala 98:55 ALU.scala 99:14]
  wire [3:0] _GEN_26 = ~opcode_4 & ~opcode_3 ? _gate_a_T : _GEN_22; // @[ALU.scala 93:49 ALU.scala 94:14]
  wire  _T_38 = ~opcode_5; // @[ALU.scala 114:66]
  wire [3:0] _GEN_30 = _T_34 ? io_in_a : snapshot_a; // @[ALU.scala 125:55 ALU.scala 126:14 ALU.scala 131:14]
  wire [3:0] _GEN_34 = _T_31 ? snapshot_a : _GEN_30; // @[ALU.scala 120:55 ALU.scala 121:14]
  wire [3:0] _GEN_38 = _T_28 ? io_in_a : _GEN_34; // @[ALU.scala 115:49 ALU.scala 116:14]
  wire [3:0] _GEN_54 = opcode_8 & opcode_6 & ~opcode_5 ? _GEN_38 : _GEN_38; // @[ALU.scala 114:74]
  wire [3:0] gate_a = opcode_8 & ~opcode_6 & opcode_5 ? _GEN_26 : _GEN_54; // @[ALU.scala 92:68]
  wire [3:0] _GEN_23 = opcode_4 & _T_27 ? io_in_b : snapshot_b; // @[ALU.scala 98:55 ALU.scala 100:14]
  wire [3:0] _GEN_27 = ~opcode_4 & ~opcode_3 ? io_in_b : _GEN_23; // @[ALU.scala 93:49 ALU.scala 95:14]
  wire [3:0] _gate_b_T = ~io_in_b; // @[ALU.scala 117:17]
  wire [3:0] _gate_b_T_2 = ~snapshot_b; // @[ALU.scala 127:17]
  wire [3:0] _GEN_31 = _T_34 ? _gate_b_T_2 : _gate_b_T_2; // @[ALU.scala 125:55 ALU.scala 127:14 ALU.scala 132:14]
  wire [3:0] _GEN_35 = _T_31 ? _gate_b_T : _GEN_31; // @[ALU.scala 120:55 ALU.scala 122:14]
  wire [3:0] _GEN_39 = _T_28 ? _gate_b_T : _GEN_35; // @[ALU.scala 115:49 ALU.scala 117:14]
  wire [3:0] _GEN_55 = opcode_8 & opcode_6 & ~opcode_5 ? _GEN_39 : _GEN_27; // @[ALU.scala 114:74]
  wire [3:0] gate_b = opcode_8 & ~opcode_6 & opcode_5 ? _GEN_27 : _GEN_55; // @[ALU.scala 92:68]
  wire [3:0] _temp_result_a_T = gate_a & gate_b; // @[ALU.scala 53:33]
  wire [3:0] _temp_result_a_T_1 = ~_temp_result_a_T; // @[ALU.scala 53:24]
  wire [3:0] _temp_result_a_T_3 = gate_a | gate_b; // @[ALU.scala 61:33]
  wire [3:0] _temp_result_a_T_4 = ~_temp_result_a_T_3; // @[ALU.scala 61:24]
  wire  _T_12 = ~opcode_8; // @[ALU.scala 67:24]
  wire [3:0] _temp_result_a_T_6 = gate_a ^ gate_b; // @[ALU.scala 69:33]
  wire [3:0] _temp_result_a_T_7 = ~_temp_result_a_T_6; // @[ALU.scala 69:24]
  wire [3:0] _GEN_4 = opcode_5 ? _temp_result_a_T_7 : _temp_result_a_T_6; // @[ALU.scala 68:28 ALU.scala 69:21 ALU.scala 72:21]
  wire  _T_18 = _T_12 & _T_1; // @[ALU.scala 75:32]
  wire [3:0] _temp_result_a_T_9 = ~gate_a; // @[ALU.scala 80:24]
  wire [3:0] _GEN_6 = opcode_5 ? _temp_result_a_T_9 : temp_result_a; // @[ALU.scala 79:34 ALU.scala 80:21 ALU.scala 33:30]
  wire [3:0] _GEN_7 = opcode_5 ? gate_b : temp_result_b; // @[ALU.scala 79:34 ALU.scala 81:21 ALU.scala 34:30]
  wire [3:0] _GEN_8 = _T_38 ? gate_a : _GEN_6; // @[ALU.scala 76:28 ALU.scala 77:21]
  wire [3:0] _GEN_9 = _T_38 ? gate_b : _GEN_7; // @[ALU.scala 76:28 ALU.scala 78:21]
  wire [3:0] _GEN_10 = _T_12 & _T_1 ? _GEN_8 : temp_result_a; // @[ALU.scala 75:53 ALU.scala 33:30]
  wire [3:0] _GEN_11 = _T_12 & _T_1 ? _GEN_9 : temp_result_b; // @[ALU.scala 75:53 ALU.scala 34:30]
  wire  _GEN_20 = _T_26 & opcode_3 ? io_validin_a : snapshot_valid_a; // @[ALU.scala 103:55 ALU.scala 106:20 ALU.scala 111:20]
  wire  _GEN_24 = opcode_4 & _T_27 ? snapshot_valid_a : _GEN_20; // @[ALU.scala 98:55 ALU.scala 101:20]
  wire  _GEN_25 = opcode_4 & _T_27 ? io_validin_b : snapshot_valid_b; // @[ALU.scala 98:55 ALU.scala 102:20]
  wire  _GEN_28 = ~opcode_4 & ~opcode_3 ? io_validin_a : _GEN_24; // @[ALU.scala 93:49 ALU.scala 96:20]
  wire  _GEN_29 = ~opcode_4 & ~opcode_3 ? io_validin_b : _GEN_25; // @[ALU.scala 93:49 ALU.scala 97:20]
  wire  _GEN_56 = opcode_8 & opcode_6 & ~opcode_5 ? _GEN_28 : _GEN_28; // @[ALU.scala 114:74]
  wire  _GEN_57 = opcode_8 & opcode_6 & ~opcode_5 ? _GEN_29 : _GEN_29; // @[ALU.scala 114:74]
  wire  gate_valid_a = opcode_8 & ~opcode_6 & opcode_5 ? _GEN_28 : _GEN_56; // @[ALU.scala 92:68]
  wire  gate_valid_b = opcode_8 & ~opcode_6 & opcode_5 ? _GEN_29 : _GEN_57; // @[ALU.scala 92:68]
  wire  _T_65 = ~opcode_0; // @[ALU.scala 178:20]
  wire  _GEN_70 = opcode_0 ? gate_valid_a : temp_valid_a; // @[ALU.scala 181:35 ALU.scala 182:20 ALU.scala 37:29]
  wire  _GEN_71 = opcode_0 ? gate_valid_b : temp_valid_b; // @[ALU.scala 181:35 ALU.scala 183:20 ALU.scala 38:29]
  assign io_out_a = temp_result_a; // @[ALU.scala 217:12]
  assign io_out_b = temp_result_b; // @[ALU.scala 218:12]
  assign io_validout_a = temp_valid_a; // @[ALU.scala 219:17]
  assign io_validout_b = temp_valid_b; // @[ALU.scala 220:17]
  always @(posedge clock) begin
    if (reset) begin // @[ALU.scala 25:27]
      snapshot_a <= 4'h0; // @[ALU.scala 25:27]
    end else if (opcode_2) begin // @[ALU.scala 160:26]
      snapshot_a <= io_in_a; // @[ALU.scala 161:16]
    end
    if (reset) begin // @[ALU.scala 26:27]
      snapshot_b <= 4'h0; // @[ALU.scala 26:27]
    end else if (opcode_1) begin // @[ALU.scala 168:26]
      snapshot_b <= io_in_b; // @[ALU.scala 169:16]
    end
    if (reset) begin // @[ALU.scala 28:33]
      snapshot_valid_a <= 1'h0; // @[ALU.scala 28:33]
    end else if (opcode_2) begin // @[ALU.scala 160:26]
      snapshot_valid_a <= io_validin_a; // @[ALU.scala 162:22]
    end
    if (reset) begin // @[ALU.scala 29:33]
      snapshot_valid_b <= 1'h0; // @[ALU.scala 29:33]
    end else if (opcode_1) begin // @[ALU.scala 168:26]
      snapshot_valid_b <= io_validin_b; // @[ALU.scala 170:22]
    end
    if (reset) begin // @[ALU.scala 33:30]
      temp_result_a <= 4'h0; // @[ALU.scala 33:30]
    end else if (opcode_8 & ~opcode_7) begin // @[ALU.scala 51:47]
      if (opcode_6 & opcode_5) begin // @[ALU.scala 52:49]
        temp_result_a <= _temp_result_a_T_1; // @[ALU.scala 53:21]
      end else begin
        temp_result_a <= _temp_result_a_T; // @[ALU.scala 56:21]
      end
    end else if (opcode_8 & opcode_7) begin // @[ALU.scala 59:53]
      if (_T_5) begin // @[ALU.scala 60:49]
        temp_result_a <= _temp_result_a_T_4; // @[ALU.scala 61:21]
      end else begin
        temp_result_a <= _temp_result_a_T_3; // @[ALU.scala 64:21]
      end
    end else if (~opcode_8 & opcode_7) begin // @[ALU.scala 67:53]
      temp_result_a <= _GEN_4;
    end else begin
      temp_result_a <= _GEN_10;
    end
    if (reset) begin // @[ALU.scala 34:30]
      temp_result_b <= 4'h0; // @[ALU.scala 34:30]
    end else if (opcode_8 & ~opcode_7) begin // @[ALU.scala 51:47]
      temp_result_b <= gate_b;
    end else if (opcode_8 & opcode_7) begin // @[ALU.scala 59:53]
      temp_result_b <= gate_b;
    end else if (~opcode_8 & opcode_7) begin // @[ALU.scala 67:53]
      temp_result_b <= gate_b;
    end else begin
      temp_result_b <= _GEN_11;
    end
    if (reset) begin // @[ALU.scala 37:29]
      temp_valid_a <= 1'h0; // @[ALU.scala 37:29]
    end else if (_T_18) begin // @[ALU.scala 177:47]
      if (~opcode_0) begin // @[ALU.scala 178:29]
        temp_valid_a <= gate_valid_a; // @[ALU.scala 179:20]
      end else begin
        temp_valid_a <= _GEN_70;
      end
    end else if (_T_65) begin // @[ALU.scala 186:29]
      temp_valid_a <= 1'h0; // @[ALU.scala 187:20]
    end else begin
      temp_valid_a <= _GEN_70;
    end
    if (reset) begin // @[ALU.scala 38:29]
      temp_valid_b <= 1'h0; // @[ALU.scala 38:29]
    end else if (_T_18) begin // @[ALU.scala 177:47]
      if (~opcode_0) begin // @[ALU.scala 178:29]
        temp_valid_b <= 1'h0; // @[ALU.scala 180:20]
      end else begin
        temp_valid_b <= _GEN_71;
      end
    end else if (_T_65) begin // @[ALU.scala 186:29]
      temp_valid_b <= gate_valid_b; // @[ALU.scala 188:20]
    end else begin
      temp_valid_b <= _GEN_71;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  snapshot_a = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  snapshot_b = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  snapshot_valid_a = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  snapshot_valid_b = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  temp_result_a = _RAND_4[3:0];
  _RAND_5 = {1{`RANDOM}};
  temp_result_b = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  temp_valid_a = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  temp_valid_b = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module PEcol(
  input          clock,
  input          reset,
  input  [3:0]   io_d_in_0_a,
  input          io_d_in_0_valid_a,
  input  [3:0]   io_d_in_0_b,
  input          io_d_in_0_valid_b,
  input  [3:0]   io_d_in_1_a,
  input          io_d_in_1_valid_a,
  input  [3:0]   io_d_in_1_b,
  input          io_d_in_1_valid_b,
  input  [3:0]   io_d_in_2_a,
  input          io_d_in_2_valid_a,
  input  [3:0]   io_d_in_2_b,
  input          io_d_in_2_valid_b,
  input  [3:0]   io_d_in_3_a,
  input          io_d_in_3_valid_a,
  input  [3:0]   io_d_in_3_b,
  input          io_d_in_3_valid_b,
  input  [3:0]   io_d_in_4_a,
  input          io_d_in_4_valid_a,
  input  [3:0]   io_d_in_4_b,
  input          io_d_in_4_valid_b,
  input  [3:0]   io_d_in_5_a,
  input          io_d_in_5_valid_a,
  input  [3:0]   io_d_in_5_b,
  input          io_d_in_5_valid_b,
  input  [3:0]   io_d_in_6_a,
  input          io_d_in_6_valid_a,
  input  [3:0]   io_d_in_6_b,
  input          io_d_in_6_valid_b,
  input  [3:0]   io_d_in_7_a,
  input          io_d_in_7_valid_a,
  input  [3:0]   io_d_in_7_b,
  input          io_d_in_7_valid_b,
  input  [3:0]   io_d_in_8_a,
  input          io_d_in_8_valid_a,
  input  [3:0]   io_d_in_8_b,
  input          io_d_in_8_valid_b,
  input  [3:0]   io_d_in_9_a,
  input          io_d_in_9_valid_a,
  input  [3:0]   io_d_in_9_b,
  input          io_d_in_9_valid_b,
  input  [3:0]   io_d_in_10_a,
  input          io_d_in_10_valid_a,
  input  [3:0]   io_d_in_10_b,
  input          io_d_in_10_valid_b,
  input  [3:0]   io_d_in_11_a,
  input          io_d_in_11_valid_a,
  input  [3:0]   io_d_in_11_b,
  input          io_d_in_11_valid_b,
  input  [3:0]   io_d_in_12_a,
  input          io_d_in_12_valid_a,
  input  [3:0]   io_d_in_12_b,
  input          io_d_in_12_valid_b,
  input  [3:0]   io_d_in_13_a,
  input          io_d_in_13_valid_a,
  input  [3:0]   io_d_in_13_b,
  input          io_d_in_13_valid_b,
  input  [3:0]   io_d_in_14_a,
  input          io_d_in_14_valid_a,
  input  [3:0]   io_d_in_14_b,
  input          io_d_in_14_valid_b,
  input  [3:0]   io_d_in_15_a,
  input          io_d_in_15_valid_a,
  input  [3:0]   io_d_in_15_b,
  input          io_d_in_15_valid_b,
  input  [3:0]   io_d_in_16_a,
  input          io_d_in_16_valid_a,
  input  [3:0]   io_d_in_16_b,
  input          io_d_in_16_valid_b,
  input  [3:0]   io_d_in_17_a,
  input          io_d_in_17_valid_a,
  input  [3:0]   io_d_in_17_b,
  input          io_d_in_17_valid_b,
  input  [3:0]   io_d_in_18_a,
  input          io_d_in_18_valid_a,
  input  [3:0]   io_d_in_18_b,
  input          io_d_in_18_valid_b,
  input  [3:0]   io_d_in_19_a,
  input          io_d_in_19_valid_a,
  input  [3:0]   io_d_in_19_b,
  input          io_d_in_19_valid_b,
  input  [3:0]   io_d_in_20_a,
  input          io_d_in_20_valid_a,
  input  [3:0]   io_d_in_20_b,
  input          io_d_in_20_valid_b,
  input  [3:0]   io_d_in_21_a,
  input          io_d_in_21_valid_a,
  input  [3:0]   io_d_in_21_b,
  input          io_d_in_21_valid_b,
  input  [3:0]   io_d_in_22_a,
  input          io_d_in_22_valid_a,
  input  [3:0]   io_d_in_22_b,
  input          io_d_in_22_valid_b,
  input  [3:0]   io_d_in_23_a,
  input          io_d_in_23_valid_a,
  input  [3:0]   io_d_in_23_b,
  input          io_d_in_23_valid_b,
  input  [3:0]   io_d_in_24_a,
  input          io_d_in_24_valid_a,
  input  [3:0]   io_d_in_24_b,
  input          io_d_in_24_valid_b,
  input  [3:0]   io_d_in_25_a,
  input          io_d_in_25_valid_a,
  input  [3:0]   io_d_in_25_b,
  input          io_d_in_25_valid_b,
  input  [3:0]   io_d_in_26_a,
  input          io_d_in_26_valid_a,
  input  [3:0]   io_d_in_26_b,
  input          io_d_in_26_valid_b,
  input  [3:0]   io_d_in_27_a,
  input          io_d_in_27_valid_a,
  input  [3:0]   io_d_in_27_b,
  input          io_d_in_27_valid_b,
  input  [3:0]   io_d_in_28_a,
  input          io_d_in_28_valid_a,
  input  [3:0]   io_d_in_28_b,
  input          io_d_in_28_valid_b,
  input  [3:0]   io_d_in_29_a,
  input          io_d_in_29_valid_a,
  input  [3:0]   io_d_in_29_b,
  input          io_d_in_29_valid_b,
  input  [3:0]   io_d_in_30_a,
  input          io_d_in_30_valid_a,
  input  [3:0]   io_d_in_30_b,
  input          io_d_in_30_valid_b,
  input  [3:0]   io_d_in_31_a,
  input          io_d_in_31_valid_a,
  input  [3:0]   io_d_in_31_b,
  input          io_d_in_31_valid_b,
  output [3:0]   io_d_out_0_a,
  output         io_d_out_0_valid_a,
  output [3:0]   io_d_out_0_b,
  output         io_d_out_0_valid_b,
  output [3:0]   io_d_out_1_a,
  output         io_d_out_1_valid_a,
  output [3:0]   io_d_out_1_b,
  output         io_d_out_1_valid_b,
  output [3:0]   io_d_out_2_a,
  output         io_d_out_2_valid_a,
  output [3:0]   io_d_out_2_b,
  output         io_d_out_2_valid_b,
  output [3:0]   io_d_out_3_a,
  output         io_d_out_3_valid_a,
  output [3:0]   io_d_out_3_b,
  output         io_d_out_3_valid_b,
  output [3:0]   io_d_out_4_a,
  output         io_d_out_4_valid_a,
  output [3:0]   io_d_out_4_b,
  output         io_d_out_4_valid_b,
  output [3:0]   io_d_out_5_a,
  output         io_d_out_5_valid_a,
  output [3:0]   io_d_out_5_b,
  output         io_d_out_5_valid_b,
  output [3:0]   io_d_out_6_a,
  output         io_d_out_6_valid_a,
  output [3:0]   io_d_out_6_b,
  output         io_d_out_6_valid_b,
  output [3:0]   io_d_out_7_a,
  output         io_d_out_7_valid_a,
  output [3:0]   io_d_out_7_b,
  output         io_d_out_7_valid_b,
  output [3:0]   io_d_out_8_a,
  output         io_d_out_8_valid_a,
  output [3:0]   io_d_out_8_b,
  output         io_d_out_8_valid_b,
  output [3:0]   io_d_out_9_a,
  output         io_d_out_9_valid_a,
  output [3:0]   io_d_out_9_b,
  output         io_d_out_9_valid_b,
  output [3:0]   io_d_out_10_a,
  output         io_d_out_10_valid_a,
  output [3:0]   io_d_out_10_b,
  output         io_d_out_10_valid_b,
  output [3:0]   io_d_out_11_a,
  output         io_d_out_11_valid_a,
  output [3:0]   io_d_out_11_b,
  output         io_d_out_11_valid_b,
  output [3:0]   io_d_out_12_a,
  output         io_d_out_12_valid_a,
  output [3:0]   io_d_out_12_b,
  output         io_d_out_12_valid_b,
  output [3:0]   io_d_out_13_a,
  output         io_d_out_13_valid_a,
  output [3:0]   io_d_out_13_b,
  output         io_d_out_13_valid_b,
  output [3:0]   io_d_out_14_a,
  output         io_d_out_14_valid_a,
  output [3:0]   io_d_out_14_b,
  output         io_d_out_14_valid_b,
  output [3:0]   io_d_out_15_a,
  output         io_d_out_15_valid_a,
  output [3:0]   io_d_out_15_b,
  output         io_d_out_15_valid_b,
  output [3:0]   io_d_out_16_a,
  output         io_d_out_16_valid_a,
  output [3:0]   io_d_out_16_b,
  output         io_d_out_16_valid_b,
  output [3:0]   io_d_out_17_a,
  output         io_d_out_17_valid_a,
  output [3:0]   io_d_out_17_b,
  output         io_d_out_17_valid_b,
  output [3:0]   io_d_out_18_a,
  output         io_d_out_18_valid_a,
  output [3:0]   io_d_out_18_b,
  output         io_d_out_18_valid_b,
  output [3:0]   io_d_out_19_a,
  output         io_d_out_19_valid_a,
  output [3:0]   io_d_out_19_b,
  output         io_d_out_19_valid_b,
  output [3:0]   io_d_out_20_a,
  output         io_d_out_20_valid_a,
  output [3:0]   io_d_out_20_b,
  output         io_d_out_20_valid_b,
  output [3:0]   io_d_out_21_a,
  output         io_d_out_21_valid_a,
  output [3:0]   io_d_out_21_b,
  output         io_d_out_21_valid_b,
  output [3:0]   io_d_out_22_a,
  output         io_d_out_22_valid_a,
  output [3:0]   io_d_out_22_b,
  output         io_d_out_22_valid_b,
  output [3:0]   io_d_out_23_a,
  output         io_d_out_23_valid_a,
  output [3:0]   io_d_out_23_b,
  output         io_d_out_23_valid_b,
  output [3:0]   io_d_out_24_a,
  output         io_d_out_24_valid_a,
  output [3:0]   io_d_out_24_b,
  output         io_d_out_24_valid_b,
  output [3:0]   io_d_out_25_a,
  output         io_d_out_25_valid_a,
  output [3:0]   io_d_out_25_b,
  output         io_d_out_25_valid_b,
  output [3:0]   io_d_out_26_a,
  output         io_d_out_26_valid_a,
  output [3:0]   io_d_out_26_b,
  output         io_d_out_26_valid_b,
  output [3:0]   io_d_out_27_a,
  output         io_d_out_27_valid_a,
  output [3:0]   io_d_out_27_b,
  output         io_d_out_27_valid_b,
  output [3:0]   io_d_out_28_a,
  output         io_d_out_28_valid_a,
  output [3:0]   io_d_out_28_b,
  output         io_d_out_28_valid_b,
  output [3:0]   io_d_out_29_a,
  output         io_d_out_29_valid_a,
  output [3:0]   io_d_out_29_b,
  output         io_d_out_29_valid_b,
  output [3:0]   io_d_out_30_a,
  output         io_d_out_30_valid_a,
  output [3:0]   io_d_out_30_b,
  output         io_d_out_30_valid_b,
  output [3:0]   io_d_out_31_a,
  output         io_d_out_31_valid_a,
  output [3:0]   io_d_out_31_b,
  output         io_d_out_31_valid_b,
  input  [7:0]   io_addrin,
  output [7:0]   io_addrout,
  input  [287:0] io_instr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  ALU64_32_0_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_0_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_0_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_0_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_0_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_0_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_0_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_0_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_0_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_0_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_0_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_1_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_1_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_1_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_1_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_1_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_1_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_1_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_1_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_1_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_1_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_1_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_2_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_2_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_2_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_2_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_2_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_2_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_2_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_2_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_2_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_2_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_2_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_3_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_3_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_3_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_3_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_3_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_3_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_3_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_3_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_3_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_3_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_3_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_4_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_4_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_4_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_4_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_4_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_4_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_4_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_4_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_4_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_4_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_4_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_5_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_5_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_5_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_5_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_5_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_5_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_5_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_5_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_5_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_5_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_5_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_6_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_6_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_6_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_6_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_6_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_6_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_6_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_6_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_6_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_6_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_6_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_7_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_7_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_7_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_7_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_7_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_7_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_7_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_7_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_7_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_7_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_7_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_8_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_8_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_8_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_8_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_8_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_8_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_8_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_8_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_8_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_8_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_8_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_9_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_9_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_9_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_9_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_9_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_9_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_9_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_9_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_9_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_9_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_9_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_10_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_10_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_10_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_10_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_10_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_10_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_10_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_10_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_10_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_10_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_10_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_11_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_11_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_11_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_11_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_11_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_11_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_11_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_11_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_11_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_11_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_11_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_12_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_12_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_12_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_12_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_12_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_12_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_12_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_12_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_12_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_12_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_12_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_13_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_13_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_13_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_13_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_13_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_13_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_13_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_13_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_13_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_13_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_13_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_14_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_14_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_14_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_14_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_14_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_14_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_14_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_14_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_14_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_14_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_14_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_15_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_15_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_15_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_15_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_15_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_15_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_15_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_15_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_15_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_15_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_15_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_16_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_16_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_16_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_16_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_16_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_16_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_16_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_16_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_16_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_16_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_16_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_17_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_17_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_17_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_17_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_17_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_17_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_17_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_17_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_17_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_17_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_17_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_18_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_18_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_18_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_18_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_18_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_18_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_18_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_18_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_18_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_18_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_18_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_19_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_19_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_19_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_19_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_19_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_19_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_19_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_19_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_19_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_19_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_19_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_20_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_20_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_20_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_20_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_20_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_20_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_20_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_20_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_20_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_20_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_20_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_21_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_21_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_21_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_21_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_21_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_21_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_21_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_21_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_21_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_21_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_21_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_22_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_22_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_22_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_22_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_22_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_22_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_22_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_22_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_22_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_22_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_22_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_23_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_23_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_23_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_23_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_23_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_23_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_23_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_23_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_23_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_23_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_23_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_24_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_24_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_24_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_24_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_24_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_24_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_24_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_24_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_24_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_24_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_24_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_25_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_25_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_25_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_25_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_25_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_25_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_25_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_25_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_25_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_25_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_25_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_26_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_26_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_26_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_26_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_26_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_26_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_26_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_26_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_26_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_26_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_26_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_27_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_27_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_27_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_27_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_27_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_27_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_27_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_27_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_27_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_27_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_27_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_28_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_28_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_28_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_28_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_28_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_28_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_28_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_28_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_28_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_28_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_28_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_29_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_29_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_29_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_29_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_29_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_29_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_29_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_29_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_29_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_29_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_29_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_30_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_30_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_30_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_30_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_30_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_30_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_30_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_30_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_30_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_30_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_30_io_validout_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_31_clock; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_31_reset; // @[BuildingBlock.scala 230:52]
  wire [8:0] ALU64_32_31_io_opcode; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_31_io_in_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_31_io_in_b; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_31_io_out_a; // @[BuildingBlock.scala 230:52]
  wire [3:0] ALU64_32_31_io_out_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_31_io_validin_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_31_io_validin_b; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_31_io_validout_a; // @[BuildingBlock.scala 230:52]
  wire  ALU64_32_31_io_validout_b; // @[BuildingBlock.scala 230:52]
  reg [7:0] addr; // @[BuildingBlock.scala 234:21]
  ALU ALU64_32_0 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_0_clock),
    .reset(ALU64_32_0_reset),
    .io_opcode(ALU64_32_0_io_opcode),
    .io_in_a(ALU64_32_0_io_in_a),
    .io_in_b(ALU64_32_0_io_in_b),
    .io_out_a(ALU64_32_0_io_out_a),
    .io_out_b(ALU64_32_0_io_out_b),
    .io_validin_a(ALU64_32_0_io_validin_a),
    .io_validin_b(ALU64_32_0_io_validin_b),
    .io_validout_a(ALU64_32_0_io_validout_a),
    .io_validout_b(ALU64_32_0_io_validout_b)
  );
  ALU ALU64_32_1 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_1_clock),
    .reset(ALU64_32_1_reset),
    .io_opcode(ALU64_32_1_io_opcode),
    .io_in_a(ALU64_32_1_io_in_a),
    .io_in_b(ALU64_32_1_io_in_b),
    .io_out_a(ALU64_32_1_io_out_a),
    .io_out_b(ALU64_32_1_io_out_b),
    .io_validin_a(ALU64_32_1_io_validin_a),
    .io_validin_b(ALU64_32_1_io_validin_b),
    .io_validout_a(ALU64_32_1_io_validout_a),
    .io_validout_b(ALU64_32_1_io_validout_b)
  );
  ALU ALU64_32_2 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_2_clock),
    .reset(ALU64_32_2_reset),
    .io_opcode(ALU64_32_2_io_opcode),
    .io_in_a(ALU64_32_2_io_in_a),
    .io_in_b(ALU64_32_2_io_in_b),
    .io_out_a(ALU64_32_2_io_out_a),
    .io_out_b(ALU64_32_2_io_out_b),
    .io_validin_a(ALU64_32_2_io_validin_a),
    .io_validin_b(ALU64_32_2_io_validin_b),
    .io_validout_a(ALU64_32_2_io_validout_a),
    .io_validout_b(ALU64_32_2_io_validout_b)
  );
  ALU ALU64_32_3 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_3_clock),
    .reset(ALU64_32_3_reset),
    .io_opcode(ALU64_32_3_io_opcode),
    .io_in_a(ALU64_32_3_io_in_a),
    .io_in_b(ALU64_32_3_io_in_b),
    .io_out_a(ALU64_32_3_io_out_a),
    .io_out_b(ALU64_32_3_io_out_b),
    .io_validin_a(ALU64_32_3_io_validin_a),
    .io_validin_b(ALU64_32_3_io_validin_b),
    .io_validout_a(ALU64_32_3_io_validout_a),
    .io_validout_b(ALU64_32_3_io_validout_b)
  );
  ALU ALU64_32_4 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_4_clock),
    .reset(ALU64_32_4_reset),
    .io_opcode(ALU64_32_4_io_opcode),
    .io_in_a(ALU64_32_4_io_in_a),
    .io_in_b(ALU64_32_4_io_in_b),
    .io_out_a(ALU64_32_4_io_out_a),
    .io_out_b(ALU64_32_4_io_out_b),
    .io_validin_a(ALU64_32_4_io_validin_a),
    .io_validin_b(ALU64_32_4_io_validin_b),
    .io_validout_a(ALU64_32_4_io_validout_a),
    .io_validout_b(ALU64_32_4_io_validout_b)
  );
  ALU ALU64_32_5 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_5_clock),
    .reset(ALU64_32_5_reset),
    .io_opcode(ALU64_32_5_io_opcode),
    .io_in_a(ALU64_32_5_io_in_a),
    .io_in_b(ALU64_32_5_io_in_b),
    .io_out_a(ALU64_32_5_io_out_a),
    .io_out_b(ALU64_32_5_io_out_b),
    .io_validin_a(ALU64_32_5_io_validin_a),
    .io_validin_b(ALU64_32_5_io_validin_b),
    .io_validout_a(ALU64_32_5_io_validout_a),
    .io_validout_b(ALU64_32_5_io_validout_b)
  );
  ALU ALU64_32_6 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_6_clock),
    .reset(ALU64_32_6_reset),
    .io_opcode(ALU64_32_6_io_opcode),
    .io_in_a(ALU64_32_6_io_in_a),
    .io_in_b(ALU64_32_6_io_in_b),
    .io_out_a(ALU64_32_6_io_out_a),
    .io_out_b(ALU64_32_6_io_out_b),
    .io_validin_a(ALU64_32_6_io_validin_a),
    .io_validin_b(ALU64_32_6_io_validin_b),
    .io_validout_a(ALU64_32_6_io_validout_a),
    .io_validout_b(ALU64_32_6_io_validout_b)
  );
  ALU ALU64_32_7 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_7_clock),
    .reset(ALU64_32_7_reset),
    .io_opcode(ALU64_32_7_io_opcode),
    .io_in_a(ALU64_32_7_io_in_a),
    .io_in_b(ALU64_32_7_io_in_b),
    .io_out_a(ALU64_32_7_io_out_a),
    .io_out_b(ALU64_32_7_io_out_b),
    .io_validin_a(ALU64_32_7_io_validin_a),
    .io_validin_b(ALU64_32_7_io_validin_b),
    .io_validout_a(ALU64_32_7_io_validout_a),
    .io_validout_b(ALU64_32_7_io_validout_b)
  );
  ALU ALU64_32_8 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_8_clock),
    .reset(ALU64_32_8_reset),
    .io_opcode(ALU64_32_8_io_opcode),
    .io_in_a(ALU64_32_8_io_in_a),
    .io_in_b(ALU64_32_8_io_in_b),
    .io_out_a(ALU64_32_8_io_out_a),
    .io_out_b(ALU64_32_8_io_out_b),
    .io_validin_a(ALU64_32_8_io_validin_a),
    .io_validin_b(ALU64_32_8_io_validin_b),
    .io_validout_a(ALU64_32_8_io_validout_a),
    .io_validout_b(ALU64_32_8_io_validout_b)
  );
  ALU ALU64_32_9 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_9_clock),
    .reset(ALU64_32_9_reset),
    .io_opcode(ALU64_32_9_io_opcode),
    .io_in_a(ALU64_32_9_io_in_a),
    .io_in_b(ALU64_32_9_io_in_b),
    .io_out_a(ALU64_32_9_io_out_a),
    .io_out_b(ALU64_32_9_io_out_b),
    .io_validin_a(ALU64_32_9_io_validin_a),
    .io_validin_b(ALU64_32_9_io_validin_b),
    .io_validout_a(ALU64_32_9_io_validout_a),
    .io_validout_b(ALU64_32_9_io_validout_b)
  );
  ALU ALU64_32_10 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_10_clock),
    .reset(ALU64_32_10_reset),
    .io_opcode(ALU64_32_10_io_opcode),
    .io_in_a(ALU64_32_10_io_in_a),
    .io_in_b(ALU64_32_10_io_in_b),
    .io_out_a(ALU64_32_10_io_out_a),
    .io_out_b(ALU64_32_10_io_out_b),
    .io_validin_a(ALU64_32_10_io_validin_a),
    .io_validin_b(ALU64_32_10_io_validin_b),
    .io_validout_a(ALU64_32_10_io_validout_a),
    .io_validout_b(ALU64_32_10_io_validout_b)
  );
  ALU ALU64_32_11 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_11_clock),
    .reset(ALU64_32_11_reset),
    .io_opcode(ALU64_32_11_io_opcode),
    .io_in_a(ALU64_32_11_io_in_a),
    .io_in_b(ALU64_32_11_io_in_b),
    .io_out_a(ALU64_32_11_io_out_a),
    .io_out_b(ALU64_32_11_io_out_b),
    .io_validin_a(ALU64_32_11_io_validin_a),
    .io_validin_b(ALU64_32_11_io_validin_b),
    .io_validout_a(ALU64_32_11_io_validout_a),
    .io_validout_b(ALU64_32_11_io_validout_b)
  );
  ALU ALU64_32_12 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_12_clock),
    .reset(ALU64_32_12_reset),
    .io_opcode(ALU64_32_12_io_opcode),
    .io_in_a(ALU64_32_12_io_in_a),
    .io_in_b(ALU64_32_12_io_in_b),
    .io_out_a(ALU64_32_12_io_out_a),
    .io_out_b(ALU64_32_12_io_out_b),
    .io_validin_a(ALU64_32_12_io_validin_a),
    .io_validin_b(ALU64_32_12_io_validin_b),
    .io_validout_a(ALU64_32_12_io_validout_a),
    .io_validout_b(ALU64_32_12_io_validout_b)
  );
  ALU ALU64_32_13 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_13_clock),
    .reset(ALU64_32_13_reset),
    .io_opcode(ALU64_32_13_io_opcode),
    .io_in_a(ALU64_32_13_io_in_a),
    .io_in_b(ALU64_32_13_io_in_b),
    .io_out_a(ALU64_32_13_io_out_a),
    .io_out_b(ALU64_32_13_io_out_b),
    .io_validin_a(ALU64_32_13_io_validin_a),
    .io_validin_b(ALU64_32_13_io_validin_b),
    .io_validout_a(ALU64_32_13_io_validout_a),
    .io_validout_b(ALU64_32_13_io_validout_b)
  );
  ALU ALU64_32_14 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_14_clock),
    .reset(ALU64_32_14_reset),
    .io_opcode(ALU64_32_14_io_opcode),
    .io_in_a(ALU64_32_14_io_in_a),
    .io_in_b(ALU64_32_14_io_in_b),
    .io_out_a(ALU64_32_14_io_out_a),
    .io_out_b(ALU64_32_14_io_out_b),
    .io_validin_a(ALU64_32_14_io_validin_a),
    .io_validin_b(ALU64_32_14_io_validin_b),
    .io_validout_a(ALU64_32_14_io_validout_a),
    .io_validout_b(ALU64_32_14_io_validout_b)
  );
  ALU ALU64_32_15 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_15_clock),
    .reset(ALU64_32_15_reset),
    .io_opcode(ALU64_32_15_io_opcode),
    .io_in_a(ALU64_32_15_io_in_a),
    .io_in_b(ALU64_32_15_io_in_b),
    .io_out_a(ALU64_32_15_io_out_a),
    .io_out_b(ALU64_32_15_io_out_b),
    .io_validin_a(ALU64_32_15_io_validin_a),
    .io_validin_b(ALU64_32_15_io_validin_b),
    .io_validout_a(ALU64_32_15_io_validout_a),
    .io_validout_b(ALU64_32_15_io_validout_b)
  );
  ALU ALU64_32_16 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_16_clock),
    .reset(ALU64_32_16_reset),
    .io_opcode(ALU64_32_16_io_opcode),
    .io_in_a(ALU64_32_16_io_in_a),
    .io_in_b(ALU64_32_16_io_in_b),
    .io_out_a(ALU64_32_16_io_out_a),
    .io_out_b(ALU64_32_16_io_out_b),
    .io_validin_a(ALU64_32_16_io_validin_a),
    .io_validin_b(ALU64_32_16_io_validin_b),
    .io_validout_a(ALU64_32_16_io_validout_a),
    .io_validout_b(ALU64_32_16_io_validout_b)
  );
  ALU ALU64_32_17 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_17_clock),
    .reset(ALU64_32_17_reset),
    .io_opcode(ALU64_32_17_io_opcode),
    .io_in_a(ALU64_32_17_io_in_a),
    .io_in_b(ALU64_32_17_io_in_b),
    .io_out_a(ALU64_32_17_io_out_a),
    .io_out_b(ALU64_32_17_io_out_b),
    .io_validin_a(ALU64_32_17_io_validin_a),
    .io_validin_b(ALU64_32_17_io_validin_b),
    .io_validout_a(ALU64_32_17_io_validout_a),
    .io_validout_b(ALU64_32_17_io_validout_b)
  );
  ALU ALU64_32_18 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_18_clock),
    .reset(ALU64_32_18_reset),
    .io_opcode(ALU64_32_18_io_opcode),
    .io_in_a(ALU64_32_18_io_in_a),
    .io_in_b(ALU64_32_18_io_in_b),
    .io_out_a(ALU64_32_18_io_out_a),
    .io_out_b(ALU64_32_18_io_out_b),
    .io_validin_a(ALU64_32_18_io_validin_a),
    .io_validin_b(ALU64_32_18_io_validin_b),
    .io_validout_a(ALU64_32_18_io_validout_a),
    .io_validout_b(ALU64_32_18_io_validout_b)
  );
  ALU ALU64_32_19 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_19_clock),
    .reset(ALU64_32_19_reset),
    .io_opcode(ALU64_32_19_io_opcode),
    .io_in_a(ALU64_32_19_io_in_a),
    .io_in_b(ALU64_32_19_io_in_b),
    .io_out_a(ALU64_32_19_io_out_a),
    .io_out_b(ALU64_32_19_io_out_b),
    .io_validin_a(ALU64_32_19_io_validin_a),
    .io_validin_b(ALU64_32_19_io_validin_b),
    .io_validout_a(ALU64_32_19_io_validout_a),
    .io_validout_b(ALU64_32_19_io_validout_b)
  );
  ALU ALU64_32_20 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_20_clock),
    .reset(ALU64_32_20_reset),
    .io_opcode(ALU64_32_20_io_opcode),
    .io_in_a(ALU64_32_20_io_in_a),
    .io_in_b(ALU64_32_20_io_in_b),
    .io_out_a(ALU64_32_20_io_out_a),
    .io_out_b(ALU64_32_20_io_out_b),
    .io_validin_a(ALU64_32_20_io_validin_a),
    .io_validin_b(ALU64_32_20_io_validin_b),
    .io_validout_a(ALU64_32_20_io_validout_a),
    .io_validout_b(ALU64_32_20_io_validout_b)
  );
  ALU ALU64_32_21 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_21_clock),
    .reset(ALU64_32_21_reset),
    .io_opcode(ALU64_32_21_io_opcode),
    .io_in_a(ALU64_32_21_io_in_a),
    .io_in_b(ALU64_32_21_io_in_b),
    .io_out_a(ALU64_32_21_io_out_a),
    .io_out_b(ALU64_32_21_io_out_b),
    .io_validin_a(ALU64_32_21_io_validin_a),
    .io_validin_b(ALU64_32_21_io_validin_b),
    .io_validout_a(ALU64_32_21_io_validout_a),
    .io_validout_b(ALU64_32_21_io_validout_b)
  );
  ALU ALU64_32_22 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_22_clock),
    .reset(ALU64_32_22_reset),
    .io_opcode(ALU64_32_22_io_opcode),
    .io_in_a(ALU64_32_22_io_in_a),
    .io_in_b(ALU64_32_22_io_in_b),
    .io_out_a(ALU64_32_22_io_out_a),
    .io_out_b(ALU64_32_22_io_out_b),
    .io_validin_a(ALU64_32_22_io_validin_a),
    .io_validin_b(ALU64_32_22_io_validin_b),
    .io_validout_a(ALU64_32_22_io_validout_a),
    .io_validout_b(ALU64_32_22_io_validout_b)
  );
  ALU ALU64_32_23 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_23_clock),
    .reset(ALU64_32_23_reset),
    .io_opcode(ALU64_32_23_io_opcode),
    .io_in_a(ALU64_32_23_io_in_a),
    .io_in_b(ALU64_32_23_io_in_b),
    .io_out_a(ALU64_32_23_io_out_a),
    .io_out_b(ALU64_32_23_io_out_b),
    .io_validin_a(ALU64_32_23_io_validin_a),
    .io_validin_b(ALU64_32_23_io_validin_b),
    .io_validout_a(ALU64_32_23_io_validout_a),
    .io_validout_b(ALU64_32_23_io_validout_b)
  );
  ALU ALU64_32_24 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_24_clock),
    .reset(ALU64_32_24_reset),
    .io_opcode(ALU64_32_24_io_opcode),
    .io_in_a(ALU64_32_24_io_in_a),
    .io_in_b(ALU64_32_24_io_in_b),
    .io_out_a(ALU64_32_24_io_out_a),
    .io_out_b(ALU64_32_24_io_out_b),
    .io_validin_a(ALU64_32_24_io_validin_a),
    .io_validin_b(ALU64_32_24_io_validin_b),
    .io_validout_a(ALU64_32_24_io_validout_a),
    .io_validout_b(ALU64_32_24_io_validout_b)
  );
  ALU ALU64_32_25 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_25_clock),
    .reset(ALU64_32_25_reset),
    .io_opcode(ALU64_32_25_io_opcode),
    .io_in_a(ALU64_32_25_io_in_a),
    .io_in_b(ALU64_32_25_io_in_b),
    .io_out_a(ALU64_32_25_io_out_a),
    .io_out_b(ALU64_32_25_io_out_b),
    .io_validin_a(ALU64_32_25_io_validin_a),
    .io_validin_b(ALU64_32_25_io_validin_b),
    .io_validout_a(ALU64_32_25_io_validout_a),
    .io_validout_b(ALU64_32_25_io_validout_b)
  );
  ALU ALU64_32_26 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_26_clock),
    .reset(ALU64_32_26_reset),
    .io_opcode(ALU64_32_26_io_opcode),
    .io_in_a(ALU64_32_26_io_in_a),
    .io_in_b(ALU64_32_26_io_in_b),
    .io_out_a(ALU64_32_26_io_out_a),
    .io_out_b(ALU64_32_26_io_out_b),
    .io_validin_a(ALU64_32_26_io_validin_a),
    .io_validin_b(ALU64_32_26_io_validin_b),
    .io_validout_a(ALU64_32_26_io_validout_a),
    .io_validout_b(ALU64_32_26_io_validout_b)
  );
  ALU ALU64_32_27 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_27_clock),
    .reset(ALU64_32_27_reset),
    .io_opcode(ALU64_32_27_io_opcode),
    .io_in_a(ALU64_32_27_io_in_a),
    .io_in_b(ALU64_32_27_io_in_b),
    .io_out_a(ALU64_32_27_io_out_a),
    .io_out_b(ALU64_32_27_io_out_b),
    .io_validin_a(ALU64_32_27_io_validin_a),
    .io_validin_b(ALU64_32_27_io_validin_b),
    .io_validout_a(ALU64_32_27_io_validout_a),
    .io_validout_b(ALU64_32_27_io_validout_b)
  );
  ALU ALU64_32_28 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_28_clock),
    .reset(ALU64_32_28_reset),
    .io_opcode(ALU64_32_28_io_opcode),
    .io_in_a(ALU64_32_28_io_in_a),
    .io_in_b(ALU64_32_28_io_in_b),
    .io_out_a(ALU64_32_28_io_out_a),
    .io_out_b(ALU64_32_28_io_out_b),
    .io_validin_a(ALU64_32_28_io_validin_a),
    .io_validin_b(ALU64_32_28_io_validin_b),
    .io_validout_a(ALU64_32_28_io_validout_a),
    .io_validout_b(ALU64_32_28_io_validout_b)
  );
  ALU ALU64_32_29 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_29_clock),
    .reset(ALU64_32_29_reset),
    .io_opcode(ALU64_32_29_io_opcode),
    .io_in_a(ALU64_32_29_io_in_a),
    .io_in_b(ALU64_32_29_io_in_b),
    .io_out_a(ALU64_32_29_io_out_a),
    .io_out_b(ALU64_32_29_io_out_b),
    .io_validin_a(ALU64_32_29_io_validin_a),
    .io_validin_b(ALU64_32_29_io_validin_b),
    .io_validout_a(ALU64_32_29_io_validout_a),
    .io_validout_b(ALU64_32_29_io_validout_b)
  );
  ALU ALU64_32_30 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_30_clock),
    .reset(ALU64_32_30_reset),
    .io_opcode(ALU64_32_30_io_opcode),
    .io_in_a(ALU64_32_30_io_in_a),
    .io_in_b(ALU64_32_30_io_in_b),
    .io_out_a(ALU64_32_30_io_out_a),
    .io_out_b(ALU64_32_30_io_out_b),
    .io_validin_a(ALU64_32_30_io_validin_a),
    .io_validin_b(ALU64_32_30_io_validin_b),
    .io_validout_a(ALU64_32_30_io_validout_a),
    .io_validout_b(ALU64_32_30_io_validout_b)
  );
  ALU ALU64_32_31 ( // @[BuildingBlock.scala 230:52]
    .clock(ALU64_32_31_clock),
    .reset(ALU64_32_31_reset),
    .io_opcode(ALU64_32_31_io_opcode),
    .io_in_a(ALU64_32_31_io_in_a),
    .io_in_b(ALU64_32_31_io_in_b),
    .io_out_a(ALU64_32_31_io_out_a),
    .io_out_b(ALU64_32_31_io_out_b),
    .io_validin_a(ALU64_32_31_io_validin_a),
    .io_validin_b(ALU64_32_31_io_validin_b),
    .io_validout_a(ALU64_32_31_io_validout_a),
    .io_validout_b(ALU64_32_31_io_validout_b)
  );
  assign io_d_out_0_a = ALU64_32_0_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_0_valid_a = ALU64_32_0_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_0_b = ALU64_32_0_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_0_valid_b = ALU64_32_0_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_1_a = ALU64_32_1_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_1_valid_a = ALU64_32_1_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_1_b = ALU64_32_1_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_1_valid_b = ALU64_32_1_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_2_a = ALU64_32_2_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_2_valid_a = ALU64_32_2_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_2_b = ALU64_32_2_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_2_valid_b = ALU64_32_2_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_3_a = ALU64_32_3_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_3_valid_a = ALU64_32_3_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_3_b = ALU64_32_3_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_3_valid_b = ALU64_32_3_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_4_a = ALU64_32_4_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_4_valid_a = ALU64_32_4_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_4_b = ALU64_32_4_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_4_valid_b = ALU64_32_4_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_5_a = ALU64_32_5_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_5_valid_a = ALU64_32_5_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_5_b = ALU64_32_5_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_5_valid_b = ALU64_32_5_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_6_a = ALU64_32_6_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_6_valid_a = ALU64_32_6_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_6_b = ALU64_32_6_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_6_valid_b = ALU64_32_6_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_7_a = ALU64_32_7_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_7_valid_a = ALU64_32_7_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_7_b = ALU64_32_7_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_7_valid_b = ALU64_32_7_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_8_a = ALU64_32_8_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_8_valid_a = ALU64_32_8_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_8_b = ALU64_32_8_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_8_valid_b = ALU64_32_8_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_9_a = ALU64_32_9_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_9_valid_a = ALU64_32_9_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_9_b = ALU64_32_9_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_9_valid_b = ALU64_32_9_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_10_a = ALU64_32_10_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_10_valid_a = ALU64_32_10_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_10_b = ALU64_32_10_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_10_valid_b = ALU64_32_10_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_11_a = ALU64_32_11_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_11_valid_a = ALU64_32_11_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_11_b = ALU64_32_11_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_11_valid_b = ALU64_32_11_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_12_a = ALU64_32_12_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_12_valid_a = ALU64_32_12_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_12_b = ALU64_32_12_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_12_valid_b = ALU64_32_12_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_13_a = ALU64_32_13_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_13_valid_a = ALU64_32_13_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_13_b = ALU64_32_13_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_13_valid_b = ALU64_32_13_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_14_a = ALU64_32_14_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_14_valid_a = ALU64_32_14_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_14_b = ALU64_32_14_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_14_valid_b = ALU64_32_14_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_15_a = ALU64_32_15_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_15_valid_a = ALU64_32_15_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_15_b = ALU64_32_15_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_15_valid_b = ALU64_32_15_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_16_a = ALU64_32_16_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_16_valid_a = ALU64_32_16_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_16_b = ALU64_32_16_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_16_valid_b = ALU64_32_16_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_17_a = ALU64_32_17_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_17_valid_a = ALU64_32_17_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_17_b = ALU64_32_17_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_17_valid_b = ALU64_32_17_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_18_a = ALU64_32_18_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_18_valid_a = ALU64_32_18_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_18_b = ALU64_32_18_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_18_valid_b = ALU64_32_18_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_19_a = ALU64_32_19_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_19_valid_a = ALU64_32_19_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_19_b = ALU64_32_19_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_19_valid_b = ALU64_32_19_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_20_a = ALU64_32_20_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_20_valid_a = ALU64_32_20_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_20_b = ALU64_32_20_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_20_valid_b = ALU64_32_20_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_21_a = ALU64_32_21_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_21_valid_a = ALU64_32_21_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_21_b = ALU64_32_21_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_21_valid_b = ALU64_32_21_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_22_a = ALU64_32_22_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_22_valid_a = ALU64_32_22_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_22_b = ALU64_32_22_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_22_valid_b = ALU64_32_22_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_23_a = ALU64_32_23_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_23_valid_a = ALU64_32_23_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_23_b = ALU64_32_23_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_23_valid_b = ALU64_32_23_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_24_a = ALU64_32_24_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_24_valid_a = ALU64_32_24_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_24_b = ALU64_32_24_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_24_valid_b = ALU64_32_24_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_25_a = ALU64_32_25_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_25_valid_a = ALU64_32_25_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_25_b = ALU64_32_25_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_25_valid_b = ALU64_32_25_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_26_a = ALU64_32_26_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_26_valid_a = ALU64_32_26_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_26_b = ALU64_32_26_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_26_valid_b = ALU64_32_26_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_27_a = ALU64_32_27_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_27_valid_a = ALU64_32_27_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_27_b = ALU64_32_27_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_27_valid_b = ALU64_32_27_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_28_a = ALU64_32_28_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_28_valid_a = ALU64_32_28_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_28_b = ALU64_32_28_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_28_valid_b = ALU64_32_28_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_29_a = ALU64_32_29_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_29_valid_a = ALU64_32_29_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_29_b = ALU64_32_29_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_29_valid_b = ALU64_32_29_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_30_a = ALU64_32_30_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_30_valid_a = ALU64_32_30_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_30_b = ALU64_32_30_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_30_valid_b = ALU64_32_30_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_d_out_31_a = ALU64_32_31_io_out_a; // @[BuildingBlock.scala 248:19]
  assign io_d_out_31_valid_a = ALU64_32_31_io_validout_a; // @[BuildingBlock.scala 250:25]
  assign io_d_out_31_b = ALU64_32_31_io_out_b; // @[BuildingBlock.scala 249:19]
  assign io_d_out_31_valid_b = ALU64_32_31_io_validout_b; // @[BuildingBlock.scala 251:25]
  assign io_addrout = addr; // @[BuildingBlock.scala 235:14]
  assign ALU64_32_0_clock = clock;
  assign ALU64_32_0_reset = reset;
  assign ALU64_32_0_io_opcode = io_instr[287:279]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_0_io_in_a = io_d_in_0_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_0_io_in_b = io_d_in_0_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_0_io_validin_a = io_d_in_0_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_0_io_validin_b = io_d_in_0_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_1_clock = clock;
  assign ALU64_32_1_reset = reset;
  assign ALU64_32_1_io_opcode = io_instr[278:270]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_1_io_in_a = io_d_in_1_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_1_io_in_b = io_d_in_1_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_1_io_validin_a = io_d_in_1_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_1_io_validin_b = io_d_in_1_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_2_clock = clock;
  assign ALU64_32_2_reset = reset;
  assign ALU64_32_2_io_opcode = io_instr[269:261]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_2_io_in_a = io_d_in_2_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_2_io_in_b = io_d_in_2_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_2_io_validin_a = io_d_in_2_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_2_io_validin_b = io_d_in_2_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_3_clock = clock;
  assign ALU64_32_3_reset = reset;
  assign ALU64_32_3_io_opcode = io_instr[260:252]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_3_io_in_a = io_d_in_3_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_3_io_in_b = io_d_in_3_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_3_io_validin_a = io_d_in_3_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_3_io_validin_b = io_d_in_3_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_4_clock = clock;
  assign ALU64_32_4_reset = reset;
  assign ALU64_32_4_io_opcode = io_instr[251:243]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_4_io_in_a = io_d_in_4_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_4_io_in_b = io_d_in_4_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_4_io_validin_a = io_d_in_4_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_4_io_validin_b = io_d_in_4_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_5_clock = clock;
  assign ALU64_32_5_reset = reset;
  assign ALU64_32_5_io_opcode = io_instr[242:234]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_5_io_in_a = io_d_in_5_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_5_io_in_b = io_d_in_5_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_5_io_validin_a = io_d_in_5_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_5_io_validin_b = io_d_in_5_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_6_clock = clock;
  assign ALU64_32_6_reset = reset;
  assign ALU64_32_6_io_opcode = io_instr[233:225]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_6_io_in_a = io_d_in_6_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_6_io_in_b = io_d_in_6_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_6_io_validin_a = io_d_in_6_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_6_io_validin_b = io_d_in_6_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_7_clock = clock;
  assign ALU64_32_7_reset = reset;
  assign ALU64_32_7_io_opcode = io_instr[224:216]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_7_io_in_a = io_d_in_7_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_7_io_in_b = io_d_in_7_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_7_io_validin_a = io_d_in_7_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_7_io_validin_b = io_d_in_7_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_8_clock = clock;
  assign ALU64_32_8_reset = reset;
  assign ALU64_32_8_io_opcode = io_instr[215:207]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_8_io_in_a = io_d_in_8_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_8_io_in_b = io_d_in_8_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_8_io_validin_a = io_d_in_8_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_8_io_validin_b = io_d_in_8_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_9_clock = clock;
  assign ALU64_32_9_reset = reset;
  assign ALU64_32_9_io_opcode = io_instr[206:198]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_9_io_in_a = io_d_in_9_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_9_io_in_b = io_d_in_9_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_9_io_validin_a = io_d_in_9_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_9_io_validin_b = io_d_in_9_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_10_clock = clock;
  assign ALU64_32_10_reset = reset;
  assign ALU64_32_10_io_opcode = io_instr[197:189]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_10_io_in_a = io_d_in_10_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_10_io_in_b = io_d_in_10_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_10_io_validin_a = io_d_in_10_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_10_io_validin_b = io_d_in_10_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_11_clock = clock;
  assign ALU64_32_11_reset = reset;
  assign ALU64_32_11_io_opcode = io_instr[188:180]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_11_io_in_a = io_d_in_11_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_11_io_in_b = io_d_in_11_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_11_io_validin_a = io_d_in_11_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_11_io_validin_b = io_d_in_11_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_12_clock = clock;
  assign ALU64_32_12_reset = reset;
  assign ALU64_32_12_io_opcode = io_instr[179:171]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_12_io_in_a = io_d_in_12_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_12_io_in_b = io_d_in_12_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_12_io_validin_a = io_d_in_12_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_12_io_validin_b = io_d_in_12_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_13_clock = clock;
  assign ALU64_32_13_reset = reset;
  assign ALU64_32_13_io_opcode = io_instr[170:162]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_13_io_in_a = io_d_in_13_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_13_io_in_b = io_d_in_13_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_13_io_validin_a = io_d_in_13_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_13_io_validin_b = io_d_in_13_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_14_clock = clock;
  assign ALU64_32_14_reset = reset;
  assign ALU64_32_14_io_opcode = io_instr[161:153]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_14_io_in_a = io_d_in_14_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_14_io_in_b = io_d_in_14_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_14_io_validin_a = io_d_in_14_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_14_io_validin_b = io_d_in_14_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_15_clock = clock;
  assign ALU64_32_15_reset = reset;
  assign ALU64_32_15_io_opcode = io_instr[152:144]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_15_io_in_a = io_d_in_15_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_15_io_in_b = io_d_in_15_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_15_io_validin_a = io_d_in_15_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_15_io_validin_b = io_d_in_15_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_16_clock = clock;
  assign ALU64_32_16_reset = reset;
  assign ALU64_32_16_io_opcode = io_instr[143:135]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_16_io_in_a = io_d_in_16_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_16_io_in_b = io_d_in_16_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_16_io_validin_a = io_d_in_16_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_16_io_validin_b = io_d_in_16_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_17_clock = clock;
  assign ALU64_32_17_reset = reset;
  assign ALU64_32_17_io_opcode = io_instr[134:126]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_17_io_in_a = io_d_in_17_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_17_io_in_b = io_d_in_17_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_17_io_validin_a = io_d_in_17_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_17_io_validin_b = io_d_in_17_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_18_clock = clock;
  assign ALU64_32_18_reset = reset;
  assign ALU64_32_18_io_opcode = io_instr[125:117]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_18_io_in_a = io_d_in_18_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_18_io_in_b = io_d_in_18_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_18_io_validin_a = io_d_in_18_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_18_io_validin_b = io_d_in_18_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_19_clock = clock;
  assign ALU64_32_19_reset = reset;
  assign ALU64_32_19_io_opcode = io_instr[116:108]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_19_io_in_a = io_d_in_19_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_19_io_in_b = io_d_in_19_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_19_io_validin_a = io_d_in_19_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_19_io_validin_b = io_d_in_19_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_20_clock = clock;
  assign ALU64_32_20_reset = reset;
  assign ALU64_32_20_io_opcode = io_instr[107:99]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_20_io_in_a = io_d_in_20_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_20_io_in_b = io_d_in_20_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_20_io_validin_a = io_d_in_20_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_20_io_validin_b = io_d_in_20_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_21_clock = clock;
  assign ALU64_32_21_reset = reset;
  assign ALU64_32_21_io_opcode = io_instr[98:90]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_21_io_in_a = io_d_in_21_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_21_io_in_b = io_d_in_21_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_21_io_validin_a = io_d_in_21_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_21_io_validin_b = io_d_in_21_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_22_clock = clock;
  assign ALU64_32_22_reset = reset;
  assign ALU64_32_22_io_opcode = io_instr[89:81]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_22_io_in_a = io_d_in_22_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_22_io_in_b = io_d_in_22_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_22_io_validin_a = io_d_in_22_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_22_io_validin_b = io_d_in_22_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_23_clock = clock;
  assign ALU64_32_23_reset = reset;
  assign ALU64_32_23_io_opcode = io_instr[80:72]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_23_io_in_a = io_d_in_23_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_23_io_in_b = io_d_in_23_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_23_io_validin_a = io_d_in_23_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_23_io_validin_b = io_d_in_23_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_24_clock = clock;
  assign ALU64_32_24_reset = reset;
  assign ALU64_32_24_io_opcode = io_instr[71:63]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_24_io_in_a = io_d_in_24_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_24_io_in_b = io_d_in_24_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_24_io_validin_a = io_d_in_24_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_24_io_validin_b = io_d_in_24_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_25_clock = clock;
  assign ALU64_32_25_reset = reset;
  assign ALU64_32_25_io_opcode = io_instr[62:54]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_25_io_in_a = io_d_in_25_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_25_io_in_b = io_d_in_25_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_25_io_validin_a = io_d_in_25_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_25_io_validin_b = io_d_in_25_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_26_clock = clock;
  assign ALU64_32_26_reset = reset;
  assign ALU64_32_26_io_opcode = io_instr[53:45]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_26_io_in_a = io_d_in_26_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_26_io_in_b = io_d_in_26_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_26_io_validin_a = io_d_in_26_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_26_io_validin_b = io_d_in_26_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_27_clock = clock;
  assign ALU64_32_27_reset = reset;
  assign ALU64_32_27_io_opcode = io_instr[44:36]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_27_io_in_a = io_d_in_27_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_27_io_in_b = io_d_in_27_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_27_io_validin_a = io_d_in_27_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_27_io_validin_b = io_d_in_27_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_28_clock = clock;
  assign ALU64_32_28_reset = reset;
  assign ALU64_32_28_io_opcode = io_instr[35:27]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_28_io_in_a = io_d_in_28_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_28_io_in_b = io_d_in_28_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_28_io_validin_a = io_d_in_28_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_28_io_validin_b = io_d_in_28_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_29_clock = clock;
  assign ALU64_32_29_reset = reset;
  assign ALU64_32_29_io_opcode = io_instr[26:18]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_29_io_in_a = io_d_in_29_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_29_io_in_b = io_d_in_29_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_29_io_validin_a = io_d_in_29_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_29_io_validin_b = io_d_in_29_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_30_clock = clock;
  assign ALU64_32_30_reset = reset;
  assign ALU64_32_30_io_opcode = io_instr[17:9]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_30_io_in_a = io_d_in_30_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_30_io_in_b = io_d_in_30_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_30_io_validin_a = io_d_in_30_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_30_io_validin_b = io_d_in_30_valid_b; // @[BuildingBlock.scala 243:30]
  assign ALU64_32_31_clock = clock;
  assign ALU64_32_31_reset = reset;
  assign ALU64_32_31_io_opcode = io_instr[8:0]; // @[BuildingBlock.scala 244:38]
  assign ALU64_32_31_io_in_a = io_d_in_31_a; // @[BuildingBlock.scala 240:25]
  assign ALU64_32_31_io_in_b = io_d_in_31_b; // @[BuildingBlock.scala 241:25]
  assign ALU64_32_31_io_validin_a = io_d_in_31_valid_a; // @[BuildingBlock.scala 242:30]
  assign ALU64_32_31_io_validin_b = io_d_in_31_valid_b; // @[BuildingBlock.scala 243:30]
  always @(posedge clock) begin
    addr <= io_addrin; // @[BuildingBlock.scala 234:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CrossBarCell(
  input  [4:0] io_fw_left,
  input  [4:0] io_fw_top,
  output [4:0] io_fw_bottom,
  output [4:0] io_fw_right,
  input        io_sel
);
  assign io_fw_bottom = io_sel ? io_fw_left : io_fw_top; // @[CrossBarSwitch.scala 15:17 CrossBarSwitch.scala 16:18 CrossBarSwitch.scala 18:18]
  assign io_fw_right = io_fw_left; // @[CrossBarSwitch.scala 14:15]
endmodule
module CrossBarSwitch(
  input        clock,
  input  [4:0] io_fw_left_0,
  input  [4:0] io_fw_left_1,
  input  [4:0] io_fw_left_2,
  input  [4:0] io_fw_left_3,
  output [4:0] io_fw_bottom_0,
  output [4:0] io_fw_bottom_1,
  output [4:0] io_fw_bottom_2,
  output [4:0] io_fw_bottom_3,
  input  [1:0] io_select_0,
  input  [1:0] io_select_1,
  input  [1:0] io_select_2,
  input  [1:0] io_select_3
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [4:0] cells_2d_0_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_0_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_0_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_0_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_0_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_1_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_1_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_1_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_1_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_1_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_2_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_2_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_2_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_2_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_2_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_3_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_3_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_3_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_3_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_3_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_4_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_4_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_4_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_4_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_4_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_5_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_5_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_5_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_5_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_5_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_6_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_6_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_6_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_6_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_6_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_7_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_7_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_7_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_7_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_7_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_8_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_8_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_8_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_8_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_8_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_9_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_9_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_9_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_9_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_9_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_10_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_10_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_10_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_10_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_10_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_11_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_11_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_11_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_11_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_11_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_12_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_12_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_12_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_12_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_12_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_13_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_13_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_13_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_13_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_13_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_14_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_14_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_14_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_14_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_14_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_15_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_15_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_15_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [4:0] cells_2d_15_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_15_io_sel; // @[CrossBarSwitch.scala 37:53]
  reg [4:0] fw_left_reg_0; // @[CrossBarSwitch.scala 33:28]
  reg [4:0] fw_left_reg_1; // @[CrossBarSwitch.scala 33:28]
  reg [4:0] fw_left_reg_2; // @[CrossBarSwitch.scala 33:28]
  reg [4:0] fw_left_reg_3; // @[CrossBarSwitch.scala 33:28]
  wire [3:0] select_onehot_0 = 4'h1 << io_select_0; // @[OneHot.scala 65:12]
  wire [3:0] select_onehot_1 = 4'h1 << io_select_1; // @[OneHot.scala 65:12]
  wire [3:0] select_onehot_2 = 4'h1 << io_select_2; // @[OneHot.scala 65:12]
  wire [3:0] select_onehot_3 = 4'h1 << io_select_3; // @[OneHot.scala 65:12]
  CrossBarCell cells_2d_0 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_0_io_fw_left),
    .io_fw_top(cells_2d_0_io_fw_top),
    .io_fw_bottom(cells_2d_0_io_fw_bottom),
    .io_fw_right(cells_2d_0_io_fw_right),
    .io_sel(cells_2d_0_io_sel)
  );
  CrossBarCell cells_2d_1 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_1_io_fw_left),
    .io_fw_top(cells_2d_1_io_fw_top),
    .io_fw_bottom(cells_2d_1_io_fw_bottom),
    .io_fw_right(cells_2d_1_io_fw_right),
    .io_sel(cells_2d_1_io_sel)
  );
  CrossBarCell cells_2d_2 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_2_io_fw_left),
    .io_fw_top(cells_2d_2_io_fw_top),
    .io_fw_bottom(cells_2d_2_io_fw_bottom),
    .io_fw_right(cells_2d_2_io_fw_right),
    .io_sel(cells_2d_2_io_sel)
  );
  CrossBarCell cells_2d_3 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_3_io_fw_left),
    .io_fw_top(cells_2d_3_io_fw_top),
    .io_fw_bottom(cells_2d_3_io_fw_bottom),
    .io_fw_right(cells_2d_3_io_fw_right),
    .io_sel(cells_2d_3_io_sel)
  );
  CrossBarCell cells_2d_4 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_4_io_fw_left),
    .io_fw_top(cells_2d_4_io_fw_top),
    .io_fw_bottom(cells_2d_4_io_fw_bottom),
    .io_fw_right(cells_2d_4_io_fw_right),
    .io_sel(cells_2d_4_io_sel)
  );
  CrossBarCell cells_2d_5 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_5_io_fw_left),
    .io_fw_top(cells_2d_5_io_fw_top),
    .io_fw_bottom(cells_2d_5_io_fw_bottom),
    .io_fw_right(cells_2d_5_io_fw_right),
    .io_sel(cells_2d_5_io_sel)
  );
  CrossBarCell cells_2d_6 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_6_io_fw_left),
    .io_fw_top(cells_2d_6_io_fw_top),
    .io_fw_bottom(cells_2d_6_io_fw_bottom),
    .io_fw_right(cells_2d_6_io_fw_right),
    .io_sel(cells_2d_6_io_sel)
  );
  CrossBarCell cells_2d_7 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_7_io_fw_left),
    .io_fw_top(cells_2d_7_io_fw_top),
    .io_fw_bottom(cells_2d_7_io_fw_bottom),
    .io_fw_right(cells_2d_7_io_fw_right),
    .io_sel(cells_2d_7_io_sel)
  );
  CrossBarCell cells_2d_8 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_8_io_fw_left),
    .io_fw_top(cells_2d_8_io_fw_top),
    .io_fw_bottom(cells_2d_8_io_fw_bottom),
    .io_fw_right(cells_2d_8_io_fw_right),
    .io_sel(cells_2d_8_io_sel)
  );
  CrossBarCell cells_2d_9 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_9_io_fw_left),
    .io_fw_top(cells_2d_9_io_fw_top),
    .io_fw_bottom(cells_2d_9_io_fw_bottom),
    .io_fw_right(cells_2d_9_io_fw_right),
    .io_sel(cells_2d_9_io_sel)
  );
  CrossBarCell cells_2d_10 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_10_io_fw_left),
    .io_fw_top(cells_2d_10_io_fw_top),
    .io_fw_bottom(cells_2d_10_io_fw_bottom),
    .io_fw_right(cells_2d_10_io_fw_right),
    .io_sel(cells_2d_10_io_sel)
  );
  CrossBarCell cells_2d_11 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_11_io_fw_left),
    .io_fw_top(cells_2d_11_io_fw_top),
    .io_fw_bottom(cells_2d_11_io_fw_bottom),
    .io_fw_right(cells_2d_11_io_fw_right),
    .io_sel(cells_2d_11_io_sel)
  );
  CrossBarCell cells_2d_12 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_12_io_fw_left),
    .io_fw_top(cells_2d_12_io_fw_top),
    .io_fw_bottom(cells_2d_12_io_fw_bottom),
    .io_fw_right(cells_2d_12_io_fw_right),
    .io_sel(cells_2d_12_io_sel)
  );
  CrossBarCell cells_2d_13 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_13_io_fw_left),
    .io_fw_top(cells_2d_13_io_fw_top),
    .io_fw_bottom(cells_2d_13_io_fw_bottom),
    .io_fw_right(cells_2d_13_io_fw_right),
    .io_sel(cells_2d_13_io_sel)
  );
  CrossBarCell cells_2d_14 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_14_io_fw_left),
    .io_fw_top(cells_2d_14_io_fw_top),
    .io_fw_bottom(cells_2d_14_io_fw_bottom),
    .io_fw_right(cells_2d_14_io_fw_right),
    .io_sel(cells_2d_14_io_sel)
  );
  CrossBarCell cells_2d_15 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_15_io_fw_left),
    .io_fw_top(cells_2d_15_io_fw_top),
    .io_fw_bottom(cells_2d_15_io_fw_bottom),
    .io_fw_right(cells_2d_15_io_fw_right),
    .io_sel(cells_2d_15_io_sel)
  );
  assign io_fw_bottom_0 = cells_2d_12_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_1 = cells_2d_13_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_2 = cells_2d_14_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_3 = cells_2d_15_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign cells_2d_0_io_fw_left = fw_left_reg_0; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_0_io_fw_top = 5'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_0_io_sel = select_onehot_0[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_1_io_fw_left = cells_2d_0_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_1_io_fw_top = 5'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_1_io_sel = select_onehot_1[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_2_io_fw_left = cells_2d_1_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_2_io_fw_top = 5'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_2_io_sel = select_onehot_2[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_3_io_fw_left = cells_2d_2_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_3_io_fw_top = 5'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_3_io_sel = select_onehot_3[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_4_io_fw_left = fw_left_reg_1; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_4_io_fw_top = cells_2d_0_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_4_io_sel = select_onehot_0[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_5_io_fw_left = cells_2d_4_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_5_io_fw_top = cells_2d_1_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_5_io_sel = select_onehot_1[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_6_io_fw_left = cells_2d_5_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_6_io_fw_top = cells_2d_2_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_6_io_sel = select_onehot_2[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_7_io_fw_left = cells_2d_6_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_7_io_fw_top = cells_2d_3_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_7_io_sel = select_onehot_3[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_8_io_fw_left = fw_left_reg_2; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_8_io_fw_top = cells_2d_4_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_8_io_sel = select_onehot_0[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_9_io_fw_left = cells_2d_8_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_9_io_fw_top = cells_2d_5_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_9_io_sel = select_onehot_1[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_10_io_fw_left = cells_2d_9_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_10_io_fw_top = cells_2d_6_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_10_io_sel = select_onehot_2[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_11_io_fw_left = cells_2d_10_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_11_io_fw_top = cells_2d_7_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_11_io_sel = select_onehot_3[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_12_io_fw_left = fw_left_reg_3; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_12_io_fw_top = cells_2d_8_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_12_io_sel = select_onehot_0[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_13_io_fw_left = cells_2d_12_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_13_io_fw_top = cells_2d_9_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_13_io_sel = select_onehot_1[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_14_io_fw_left = cells_2d_13_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_14_io_fw_top = cells_2d_10_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_14_io_sel = select_onehot_2[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_15_io_fw_left = cells_2d_14_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_15_io_fw_top = cells_2d_11_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_15_io_sel = select_onehot_3[3]; // @[CrossBarSwitch.scala 70:44]
  always @(posedge clock) begin
    fw_left_reg_0 <= io_fw_left_0; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_1 <= io_fw_left_1; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_2 <= io_fw_left_2; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_3 <= io_fw_left_3; // @[CrossBarSwitch.scala 33:28]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fw_left_reg_0 = _RAND_0[4:0];
  _RAND_1 = {1{`RANDOM}};
  fw_left_reg_1 = _RAND_1[4:0];
  _RAND_2 = {1{`RANDOM}};
  fw_left_reg_2 = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  fw_left_reg_3 = _RAND_3[4:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOScell4(
  input        clock,
  input  [4:0] io_in4_0,
  input  [4:0] io_in4_1,
  input  [4:0] io_in4_2,
  input  [4:0] io_in4_3,
  output [4:0] io_out4_0,
  output [4:0] io_out4_1,
  output [4:0] io_out4_2,
  output [4:0] io_out4_3,
  input  [7:0] io_ctrl
);
  wire  CrossBarSwitch_clock; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_left_0; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_left_1; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_left_2; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_left_3; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_bottom_0; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_bottom_1; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_bottom_2; // @[BuildingBlock.scala 18:21]
  wire [4:0] CrossBarSwitch_io_fw_bottom_3; // @[BuildingBlock.scala 18:21]
  wire [1:0] CrossBarSwitch_io_select_0; // @[BuildingBlock.scala 18:21]
  wire [1:0] CrossBarSwitch_io_select_1; // @[BuildingBlock.scala 18:21]
  wire [1:0] CrossBarSwitch_io_select_2; // @[BuildingBlock.scala 18:21]
  wire [1:0] CrossBarSwitch_io_select_3; // @[BuildingBlock.scala 18:21]
  CrossBarSwitch CrossBarSwitch ( // @[BuildingBlock.scala 18:21]
    .clock(CrossBarSwitch_clock),
    .io_fw_left_0(CrossBarSwitch_io_fw_left_0),
    .io_fw_left_1(CrossBarSwitch_io_fw_left_1),
    .io_fw_left_2(CrossBarSwitch_io_fw_left_2),
    .io_fw_left_3(CrossBarSwitch_io_fw_left_3),
    .io_fw_bottom_0(CrossBarSwitch_io_fw_bottom_0),
    .io_fw_bottom_1(CrossBarSwitch_io_fw_bottom_1),
    .io_fw_bottom_2(CrossBarSwitch_io_fw_bottom_2),
    .io_fw_bottom_3(CrossBarSwitch_io_fw_bottom_3),
    .io_select_0(CrossBarSwitch_io_select_0),
    .io_select_1(CrossBarSwitch_io_select_1),
    .io_select_2(CrossBarSwitch_io_select_2),
    .io_select_3(CrossBarSwitch_io_select_3)
  );
  assign io_out4_0 = CrossBarSwitch_io_fw_bottom_0; // @[BuildingBlock.scala 23:11]
  assign io_out4_1 = CrossBarSwitch_io_fw_bottom_1; // @[BuildingBlock.scala 23:11]
  assign io_out4_2 = CrossBarSwitch_io_fw_bottom_2; // @[BuildingBlock.scala 23:11]
  assign io_out4_3 = CrossBarSwitch_io_fw_bottom_3; // @[BuildingBlock.scala 23:11]
  assign CrossBarSwitch_clock = clock;
  assign CrossBarSwitch_io_fw_left_0 = io_in4_0; // @[BuildingBlock.scala 22:17]
  assign CrossBarSwitch_io_fw_left_1 = io_in4_1; // @[BuildingBlock.scala 22:17]
  assign CrossBarSwitch_io_fw_left_2 = io_in4_2; // @[BuildingBlock.scala 22:17]
  assign CrossBarSwitch_io_fw_left_3 = io_in4_3; // @[BuildingBlock.scala 22:17]
  assign CrossBarSwitch_io_select_0 = io_ctrl[7:6]; // @[BuildingBlock.scala 20:31]
  assign CrossBarSwitch_io_select_1 = io_ctrl[5:4]; // @[BuildingBlock.scala 20:31]
  assign CrossBarSwitch_io_select_2 = io_ctrl[3:2]; // @[BuildingBlock.scala 20:31]
  assign CrossBarSwitch_io_select_3 = io_ctrl[1:0]; // @[BuildingBlock.scala 20:31]
endmodule
module CLOSingress1(
  input          clock,
  input  [3:0]   io_in64_0,
  input  [3:0]   io_in64_1,
  input  [3:0]   io_in64_2,
  input  [3:0]   io_in64_3,
  input  [3:0]   io_in64_4,
  input  [3:0]   io_in64_5,
  input  [3:0]   io_in64_6,
  input  [3:0]   io_in64_7,
  input  [3:0]   io_in64_8,
  input  [3:0]   io_in64_9,
  input  [3:0]   io_in64_10,
  input  [3:0]   io_in64_11,
  input  [3:0]   io_in64_12,
  input  [3:0]   io_in64_13,
  input  [3:0]   io_in64_14,
  input  [3:0]   io_in64_15,
  input  [3:0]   io_in64_16,
  input  [3:0]   io_in64_17,
  input  [3:0]   io_in64_18,
  input  [3:0]   io_in64_19,
  input  [3:0]   io_in64_20,
  input  [3:0]   io_in64_21,
  input  [3:0]   io_in64_22,
  input  [3:0]   io_in64_23,
  input  [3:0]   io_in64_24,
  input  [3:0]   io_in64_25,
  input  [3:0]   io_in64_26,
  input  [3:0]   io_in64_27,
  input  [3:0]   io_in64_28,
  input  [3:0]   io_in64_29,
  input  [3:0]   io_in64_30,
  input  [3:0]   io_in64_31,
  input  [3:0]   io_in64_32,
  input  [3:0]   io_in64_33,
  input  [3:0]   io_in64_34,
  input  [3:0]   io_in64_35,
  input  [3:0]   io_in64_36,
  input  [3:0]   io_in64_37,
  input  [3:0]   io_in64_38,
  input  [3:0]   io_in64_39,
  input  [3:0]   io_in64_40,
  input  [3:0]   io_in64_41,
  input  [3:0]   io_in64_42,
  input  [3:0]   io_in64_43,
  input  [3:0]   io_in64_44,
  input  [3:0]   io_in64_45,
  input  [3:0]   io_in64_46,
  input  [3:0]   io_in64_47,
  input  [3:0]   io_in64_48,
  input  [3:0]   io_in64_49,
  input  [3:0]   io_in64_50,
  input  [3:0]   io_in64_51,
  input  [3:0]   io_in64_52,
  input  [3:0]   io_in64_53,
  input  [3:0]   io_in64_54,
  input  [3:0]   io_in64_55,
  input  [3:0]   io_in64_56,
  input  [3:0]   io_in64_57,
  input  [3:0]   io_in64_58,
  input  [3:0]   io_in64_59,
  input  [3:0]   io_in64_60,
  input  [3:0]   io_in64_61,
  input  [3:0]   io_in64_62,
  input  [3:0]   io_in64_63,
  input          io_validin64_0,
  input          io_validin64_1,
  input          io_validin64_2,
  input          io_validin64_3,
  input          io_validin64_4,
  input          io_validin64_5,
  input          io_validin64_6,
  input          io_validin64_7,
  input          io_validin64_8,
  input          io_validin64_9,
  input          io_validin64_10,
  input          io_validin64_11,
  input          io_validin64_12,
  input          io_validin64_13,
  input          io_validin64_14,
  input          io_validin64_15,
  input          io_validin64_16,
  input          io_validin64_17,
  input          io_validin64_18,
  input          io_validin64_19,
  input          io_validin64_20,
  input          io_validin64_21,
  input          io_validin64_22,
  input          io_validin64_23,
  input          io_validin64_24,
  input          io_validin64_25,
  input          io_validin64_26,
  input          io_validin64_27,
  input          io_validin64_28,
  input          io_validin64_29,
  input          io_validin64_30,
  input          io_validin64_31,
  input          io_validin64_32,
  input          io_validin64_33,
  input          io_validin64_34,
  input          io_validin64_35,
  input          io_validin64_36,
  input          io_validin64_37,
  input          io_validin64_38,
  input          io_validin64_39,
  input          io_validin64_40,
  input          io_validin64_41,
  input          io_validin64_42,
  input          io_validin64_43,
  input          io_validin64_44,
  input          io_validin64_45,
  input          io_validin64_46,
  input          io_validin64_47,
  input          io_validin64_48,
  input          io_validin64_49,
  input          io_validin64_50,
  input          io_validin64_51,
  input          io_validin64_52,
  input          io_validin64_53,
  input          io_validin64_54,
  input          io_validin64_55,
  input          io_validin64_56,
  input          io_validin64_57,
  input          io_validin64_58,
  input          io_validin64_59,
  input          io_validin64_60,
  input          io_validin64_61,
  input          io_validin64_62,
  input          io_validin64_63,
  input  [7:0]   io_addrin,
  output [3:0]   io_out64_0,
  output [3:0]   io_out64_1,
  output [3:0]   io_out64_2,
  output [3:0]   io_out64_3,
  output [3:0]   io_out64_4,
  output [3:0]   io_out64_5,
  output [3:0]   io_out64_6,
  output [3:0]   io_out64_7,
  output [3:0]   io_out64_8,
  output [3:0]   io_out64_9,
  output [3:0]   io_out64_10,
  output [3:0]   io_out64_11,
  output [3:0]   io_out64_12,
  output [3:0]   io_out64_13,
  output [3:0]   io_out64_14,
  output [3:0]   io_out64_15,
  output [3:0]   io_out64_16,
  output [3:0]   io_out64_17,
  output [3:0]   io_out64_18,
  output [3:0]   io_out64_19,
  output [3:0]   io_out64_20,
  output [3:0]   io_out64_21,
  output [3:0]   io_out64_22,
  output [3:0]   io_out64_23,
  output [3:0]   io_out64_24,
  output [3:0]   io_out64_25,
  output [3:0]   io_out64_26,
  output [3:0]   io_out64_27,
  output [3:0]   io_out64_28,
  output [3:0]   io_out64_29,
  output [3:0]   io_out64_30,
  output [3:0]   io_out64_31,
  output [3:0]   io_out64_32,
  output [3:0]   io_out64_33,
  output [3:0]   io_out64_34,
  output [3:0]   io_out64_35,
  output [3:0]   io_out64_36,
  output [3:0]   io_out64_37,
  output [3:0]   io_out64_38,
  output [3:0]   io_out64_39,
  output [3:0]   io_out64_40,
  output [3:0]   io_out64_41,
  output [3:0]   io_out64_42,
  output [3:0]   io_out64_43,
  output [3:0]   io_out64_44,
  output [3:0]   io_out64_45,
  output [3:0]   io_out64_46,
  output [3:0]   io_out64_47,
  output [3:0]   io_out64_48,
  output [3:0]   io_out64_49,
  output [3:0]   io_out64_50,
  output [3:0]   io_out64_51,
  output [3:0]   io_out64_52,
  output [3:0]   io_out64_53,
  output [3:0]   io_out64_54,
  output [3:0]   io_out64_55,
  output [3:0]   io_out64_56,
  output [3:0]   io_out64_57,
  output [3:0]   io_out64_58,
  output [3:0]   io_out64_59,
  output [3:0]   io_out64_60,
  output [3:0]   io_out64_61,
  output [3:0]   io_out64_62,
  output [3:0]   io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  ingress1_0_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_0_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_0_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_1_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_1_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_1_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_2_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_2_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_2_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_3_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_3_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_3_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_4_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_4_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_4_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_5_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_5_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_5_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_6_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_6_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_6_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_7_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_7_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_7_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_8_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_8_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_8_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_9_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_9_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_9_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_10_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_10_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_10_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_11_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_11_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_11_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_12_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_12_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_12_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_13_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_13_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_13_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_14_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_14_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_14_io_ctrl; // @[BuildingBlock.scala 39:52]
  wire  ingress1_15_clock; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_in4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_in4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_in4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_in4_3; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_out4_0; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_out4_1; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_out4_2; // @[BuildingBlock.scala 39:52]
  wire [4:0] ingress1_15_io_out4_3; // @[BuildingBlock.scala 39:52]
  wire [7:0] ingress1_15_io_ctrl; // @[BuildingBlock.scala 39:52]
  reg [7:0] addr; // @[BuildingBlock.scala 42:21]
  CLOScell4 ingress1_0 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_0_clock),
    .io_in4_0(ingress1_0_io_in4_0),
    .io_in4_1(ingress1_0_io_in4_1),
    .io_in4_2(ingress1_0_io_in4_2),
    .io_in4_3(ingress1_0_io_in4_3),
    .io_out4_0(ingress1_0_io_out4_0),
    .io_out4_1(ingress1_0_io_out4_1),
    .io_out4_2(ingress1_0_io_out4_2),
    .io_out4_3(ingress1_0_io_out4_3),
    .io_ctrl(ingress1_0_io_ctrl)
  );
  CLOScell4 ingress1_1 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_1_clock),
    .io_in4_0(ingress1_1_io_in4_0),
    .io_in4_1(ingress1_1_io_in4_1),
    .io_in4_2(ingress1_1_io_in4_2),
    .io_in4_3(ingress1_1_io_in4_3),
    .io_out4_0(ingress1_1_io_out4_0),
    .io_out4_1(ingress1_1_io_out4_1),
    .io_out4_2(ingress1_1_io_out4_2),
    .io_out4_3(ingress1_1_io_out4_3),
    .io_ctrl(ingress1_1_io_ctrl)
  );
  CLOScell4 ingress1_2 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_2_clock),
    .io_in4_0(ingress1_2_io_in4_0),
    .io_in4_1(ingress1_2_io_in4_1),
    .io_in4_2(ingress1_2_io_in4_2),
    .io_in4_3(ingress1_2_io_in4_3),
    .io_out4_0(ingress1_2_io_out4_0),
    .io_out4_1(ingress1_2_io_out4_1),
    .io_out4_2(ingress1_2_io_out4_2),
    .io_out4_3(ingress1_2_io_out4_3),
    .io_ctrl(ingress1_2_io_ctrl)
  );
  CLOScell4 ingress1_3 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_3_clock),
    .io_in4_0(ingress1_3_io_in4_0),
    .io_in4_1(ingress1_3_io_in4_1),
    .io_in4_2(ingress1_3_io_in4_2),
    .io_in4_3(ingress1_3_io_in4_3),
    .io_out4_0(ingress1_3_io_out4_0),
    .io_out4_1(ingress1_3_io_out4_1),
    .io_out4_2(ingress1_3_io_out4_2),
    .io_out4_3(ingress1_3_io_out4_3),
    .io_ctrl(ingress1_3_io_ctrl)
  );
  CLOScell4 ingress1_4 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_4_clock),
    .io_in4_0(ingress1_4_io_in4_0),
    .io_in4_1(ingress1_4_io_in4_1),
    .io_in4_2(ingress1_4_io_in4_2),
    .io_in4_3(ingress1_4_io_in4_3),
    .io_out4_0(ingress1_4_io_out4_0),
    .io_out4_1(ingress1_4_io_out4_1),
    .io_out4_2(ingress1_4_io_out4_2),
    .io_out4_3(ingress1_4_io_out4_3),
    .io_ctrl(ingress1_4_io_ctrl)
  );
  CLOScell4 ingress1_5 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_5_clock),
    .io_in4_0(ingress1_5_io_in4_0),
    .io_in4_1(ingress1_5_io_in4_1),
    .io_in4_2(ingress1_5_io_in4_2),
    .io_in4_3(ingress1_5_io_in4_3),
    .io_out4_0(ingress1_5_io_out4_0),
    .io_out4_1(ingress1_5_io_out4_1),
    .io_out4_2(ingress1_5_io_out4_2),
    .io_out4_3(ingress1_5_io_out4_3),
    .io_ctrl(ingress1_5_io_ctrl)
  );
  CLOScell4 ingress1_6 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_6_clock),
    .io_in4_0(ingress1_6_io_in4_0),
    .io_in4_1(ingress1_6_io_in4_1),
    .io_in4_2(ingress1_6_io_in4_2),
    .io_in4_3(ingress1_6_io_in4_3),
    .io_out4_0(ingress1_6_io_out4_0),
    .io_out4_1(ingress1_6_io_out4_1),
    .io_out4_2(ingress1_6_io_out4_2),
    .io_out4_3(ingress1_6_io_out4_3),
    .io_ctrl(ingress1_6_io_ctrl)
  );
  CLOScell4 ingress1_7 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_7_clock),
    .io_in4_0(ingress1_7_io_in4_0),
    .io_in4_1(ingress1_7_io_in4_1),
    .io_in4_2(ingress1_7_io_in4_2),
    .io_in4_3(ingress1_7_io_in4_3),
    .io_out4_0(ingress1_7_io_out4_0),
    .io_out4_1(ingress1_7_io_out4_1),
    .io_out4_2(ingress1_7_io_out4_2),
    .io_out4_3(ingress1_7_io_out4_3),
    .io_ctrl(ingress1_7_io_ctrl)
  );
  CLOScell4 ingress1_8 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_8_clock),
    .io_in4_0(ingress1_8_io_in4_0),
    .io_in4_1(ingress1_8_io_in4_1),
    .io_in4_2(ingress1_8_io_in4_2),
    .io_in4_3(ingress1_8_io_in4_3),
    .io_out4_0(ingress1_8_io_out4_0),
    .io_out4_1(ingress1_8_io_out4_1),
    .io_out4_2(ingress1_8_io_out4_2),
    .io_out4_3(ingress1_8_io_out4_3),
    .io_ctrl(ingress1_8_io_ctrl)
  );
  CLOScell4 ingress1_9 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_9_clock),
    .io_in4_0(ingress1_9_io_in4_0),
    .io_in4_1(ingress1_9_io_in4_1),
    .io_in4_2(ingress1_9_io_in4_2),
    .io_in4_3(ingress1_9_io_in4_3),
    .io_out4_0(ingress1_9_io_out4_0),
    .io_out4_1(ingress1_9_io_out4_1),
    .io_out4_2(ingress1_9_io_out4_2),
    .io_out4_3(ingress1_9_io_out4_3),
    .io_ctrl(ingress1_9_io_ctrl)
  );
  CLOScell4 ingress1_10 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_10_clock),
    .io_in4_0(ingress1_10_io_in4_0),
    .io_in4_1(ingress1_10_io_in4_1),
    .io_in4_2(ingress1_10_io_in4_2),
    .io_in4_3(ingress1_10_io_in4_3),
    .io_out4_0(ingress1_10_io_out4_0),
    .io_out4_1(ingress1_10_io_out4_1),
    .io_out4_2(ingress1_10_io_out4_2),
    .io_out4_3(ingress1_10_io_out4_3),
    .io_ctrl(ingress1_10_io_ctrl)
  );
  CLOScell4 ingress1_11 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_11_clock),
    .io_in4_0(ingress1_11_io_in4_0),
    .io_in4_1(ingress1_11_io_in4_1),
    .io_in4_2(ingress1_11_io_in4_2),
    .io_in4_3(ingress1_11_io_in4_3),
    .io_out4_0(ingress1_11_io_out4_0),
    .io_out4_1(ingress1_11_io_out4_1),
    .io_out4_2(ingress1_11_io_out4_2),
    .io_out4_3(ingress1_11_io_out4_3),
    .io_ctrl(ingress1_11_io_ctrl)
  );
  CLOScell4 ingress1_12 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_12_clock),
    .io_in4_0(ingress1_12_io_in4_0),
    .io_in4_1(ingress1_12_io_in4_1),
    .io_in4_2(ingress1_12_io_in4_2),
    .io_in4_3(ingress1_12_io_in4_3),
    .io_out4_0(ingress1_12_io_out4_0),
    .io_out4_1(ingress1_12_io_out4_1),
    .io_out4_2(ingress1_12_io_out4_2),
    .io_out4_3(ingress1_12_io_out4_3),
    .io_ctrl(ingress1_12_io_ctrl)
  );
  CLOScell4 ingress1_13 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_13_clock),
    .io_in4_0(ingress1_13_io_in4_0),
    .io_in4_1(ingress1_13_io_in4_1),
    .io_in4_2(ingress1_13_io_in4_2),
    .io_in4_3(ingress1_13_io_in4_3),
    .io_out4_0(ingress1_13_io_out4_0),
    .io_out4_1(ingress1_13_io_out4_1),
    .io_out4_2(ingress1_13_io_out4_2),
    .io_out4_3(ingress1_13_io_out4_3),
    .io_ctrl(ingress1_13_io_ctrl)
  );
  CLOScell4 ingress1_14 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_14_clock),
    .io_in4_0(ingress1_14_io_in4_0),
    .io_in4_1(ingress1_14_io_in4_1),
    .io_in4_2(ingress1_14_io_in4_2),
    .io_in4_3(ingress1_14_io_in4_3),
    .io_out4_0(ingress1_14_io_out4_0),
    .io_out4_1(ingress1_14_io_out4_1),
    .io_out4_2(ingress1_14_io_out4_2),
    .io_out4_3(ingress1_14_io_out4_3),
    .io_ctrl(ingress1_14_io_ctrl)
  );
  CLOScell4 ingress1_15 ( // @[BuildingBlock.scala 39:52]
    .clock(ingress1_15_clock),
    .io_in4_0(ingress1_15_io_in4_0),
    .io_in4_1(ingress1_15_io_in4_1),
    .io_in4_2(ingress1_15_io_in4_2),
    .io_in4_3(ingress1_15_io_in4_3),
    .io_out4_0(ingress1_15_io_out4_0),
    .io_out4_1(ingress1_15_io_out4_1),
    .io_out4_2(ingress1_15_io_out4_2),
    .io_out4_3(ingress1_15_io_out4_3),
    .io_ctrl(ingress1_15_io_ctrl)
  );
  assign io_out64_0 = ingress1_0_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_1 = ingress1_1_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_2 = ingress1_2_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_3 = ingress1_3_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_4 = ingress1_4_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_5 = ingress1_5_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_6 = ingress1_6_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_7 = ingress1_7_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_8 = ingress1_8_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_9 = ingress1_9_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_10 = ingress1_10_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_11 = ingress1_11_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_12 = ingress1_12_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_13 = ingress1_13_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_14 = ingress1_14_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_15 = ingress1_15_io_out4_0[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_16 = ingress1_0_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_17 = ingress1_1_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_18 = ingress1_2_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_19 = ingress1_3_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_20 = ingress1_4_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_21 = ingress1_5_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_22 = ingress1_6_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_23 = ingress1_7_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_24 = ingress1_8_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_25 = ingress1_9_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_26 = ingress1_10_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_27 = ingress1_11_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_28 = ingress1_12_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_29 = ingress1_13_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_30 = ingress1_14_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_31 = ingress1_15_io_out4_1[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_32 = ingress1_0_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_33 = ingress1_1_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_34 = ingress1_2_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_35 = ingress1_3_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_36 = ingress1_4_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_37 = ingress1_5_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_38 = ingress1_6_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_39 = ingress1_7_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_40 = ingress1_8_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_41 = ingress1_9_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_42 = ingress1_10_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_43 = ingress1_11_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_44 = ingress1_12_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_45 = ingress1_13_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_46 = ingress1_14_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_47 = ingress1_15_io_out4_2[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_48 = ingress1_0_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_49 = ingress1_1_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_50 = ingress1_2_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_51 = ingress1_3_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_52 = ingress1_4_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_53 = ingress1_5_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_54 = ingress1_6_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_55 = ingress1_7_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_56 = ingress1_8_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_57 = ingress1_9_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_58 = ingress1_10_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_59 = ingress1_11_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_60 = ingress1_12_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_61 = ingress1_13_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_62 = ingress1_14_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_out64_63 = ingress1_15_io_out4_3[3:0]; // @[BuildingBlock.scala 53:49]
  assign io_validout64_0 = ingress1_0_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_1 = ingress1_1_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_2 = ingress1_2_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_3 = ingress1_3_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_4 = ingress1_4_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_5 = ingress1_5_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_6 = ingress1_6_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_7 = ingress1_7_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_8 = ingress1_8_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_9 = ingress1_9_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_10 = ingress1_10_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_11 = ingress1_11_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_12 = ingress1_12_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_13 = ingress1_13_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_14 = ingress1_14_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_15 = ingress1_15_io_out4_0[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_16 = ingress1_0_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_17 = ingress1_1_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_18 = ingress1_2_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_19 = ingress1_3_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_20 = ingress1_4_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_21 = ingress1_5_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_22 = ingress1_6_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_23 = ingress1_7_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_24 = ingress1_8_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_25 = ingress1_9_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_26 = ingress1_10_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_27 = ingress1_11_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_28 = ingress1_12_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_29 = ingress1_13_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_30 = ingress1_14_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_31 = ingress1_15_io_out4_1[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_32 = ingress1_0_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_33 = ingress1_1_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_34 = ingress1_2_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_35 = ingress1_3_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_36 = ingress1_4_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_37 = ingress1_5_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_38 = ingress1_6_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_39 = ingress1_7_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_40 = ingress1_8_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_41 = ingress1_9_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_42 = ingress1_10_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_43 = ingress1_11_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_44 = ingress1_12_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_45 = ingress1_13_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_46 = ingress1_14_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_47 = ingress1_15_io_out4_2[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_48 = ingress1_0_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_49 = ingress1_1_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_50 = ingress1_2_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_51 = ingress1_3_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_52 = ingress1_4_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_53 = ingress1_5_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_54 = ingress1_6_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_55 = ingress1_7_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_56 = ingress1_8_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_57 = ingress1_9_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_58 = ingress1_10_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_59 = ingress1_11_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_60 = ingress1_12_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_61 = ingress1_13_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_62 = ingress1_14_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_validout64_63 = ingress1_15_io_out4_3[4]; // @[BuildingBlock.scala 54:54]
  assign io_addrout = addr; // @[BuildingBlock.scala 43:14]
  assign ingress1_0_clock = clock;
  assign ingress1_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign ingress1_0_io_in4_1 = {io_validin64_1,io_in64_1}; // @[Cat.scala 30:58]
  assign ingress1_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign ingress1_0_io_in4_3 = {io_validin64_3,io_in64_3}; // @[Cat.scala 30:58]
  assign ingress1_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 58:35]
  assign ingress1_1_clock = clock;
  assign ingress1_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign ingress1_1_io_in4_1 = {io_validin64_5,io_in64_5}; // @[Cat.scala 30:58]
  assign ingress1_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign ingress1_1_io_in4_3 = {io_validin64_7,io_in64_7}; // @[Cat.scala 30:58]
  assign ingress1_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 58:35]
  assign ingress1_2_clock = clock;
  assign ingress1_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign ingress1_2_io_in4_1 = {io_validin64_9,io_in64_9}; // @[Cat.scala 30:58]
  assign ingress1_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign ingress1_2_io_in4_3 = {io_validin64_11,io_in64_11}; // @[Cat.scala 30:58]
  assign ingress1_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 58:35]
  assign ingress1_3_clock = clock;
  assign ingress1_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign ingress1_3_io_in4_1 = {io_validin64_13,io_in64_13}; // @[Cat.scala 30:58]
  assign ingress1_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign ingress1_3_io_in4_3 = {io_validin64_15,io_in64_15}; // @[Cat.scala 30:58]
  assign ingress1_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 58:35]
  assign ingress1_4_clock = clock;
  assign ingress1_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign ingress1_4_io_in4_1 = {io_validin64_17,io_in64_17}; // @[Cat.scala 30:58]
  assign ingress1_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign ingress1_4_io_in4_3 = {io_validin64_19,io_in64_19}; // @[Cat.scala 30:58]
  assign ingress1_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 58:35]
  assign ingress1_5_clock = clock;
  assign ingress1_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign ingress1_5_io_in4_1 = {io_validin64_21,io_in64_21}; // @[Cat.scala 30:58]
  assign ingress1_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign ingress1_5_io_in4_3 = {io_validin64_23,io_in64_23}; // @[Cat.scala 30:58]
  assign ingress1_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 58:35]
  assign ingress1_6_clock = clock;
  assign ingress1_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign ingress1_6_io_in4_1 = {io_validin64_25,io_in64_25}; // @[Cat.scala 30:58]
  assign ingress1_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign ingress1_6_io_in4_3 = {io_validin64_27,io_in64_27}; // @[Cat.scala 30:58]
  assign ingress1_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 58:35]
  assign ingress1_7_clock = clock;
  assign ingress1_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign ingress1_7_io_in4_1 = {io_validin64_29,io_in64_29}; // @[Cat.scala 30:58]
  assign ingress1_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign ingress1_7_io_in4_3 = {io_validin64_31,io_in64_31}; // @[Cat.scala 30:58]
  assign ingress1_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 58:35]
  assign ingress1_8_clock = clock;
  assign ingress1_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign ingress1_8_io_in4_1 = {io_validin64_33,io_in64_33}; // @[Cat.scala 30:58]
  assign ingress1_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign ingress1_8_io_in4_3 = {io_validin64_35,io_in64_35}; // @[Cat.scala 30:58]
  assign ingress1_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 58:35]
  assign ingress1_9_clock = clock;
  assign ingress1_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign ingress1_9_io_in4_1 = {io_validin64_37,io_in64_37}; // @[Cat.scala 30:58]
  assign ingress1_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign ingress1_9_io_in4_3 = {io_validin64_39,io_in64_39}; // @[Cat.scala 30:58]
  assign ingress1_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 58:35]
  assign ingress1_10_clock = clock;
  assign ingress1_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign ingress1_10_io_in4_1 = {io_validin64_41,io_in64_41}; // @[Cat.scala 30:58]
  assign ingress1_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign ingress1_10_io_in4_3 = {io_validin64_43,io_in64_43}; // @[Cat.scala 30:58]
  assign ingress1_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 58:35]
  assign ingress1_11_clock = clock;
  assign ingress1_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign ingress1_11_io_in4_1 = {io_validin64_45,io_in64_45}; // @[Cat.scala 30:58]
  assign ingress1_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign ingress1_11_io_in4_3 = {io_validin64_47,io_in64_47}; // @[Cat.scala 30:58]
  assign ingress1_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 58:35]
  assign ingress1_12_clock = clock;
  assign ingress1_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign ingress1_12_io_in4_1 = {io_validin64_49,io_in64_49}; // @[Cat.scala 30:58]
  assign ingress1_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign ingress1_12_io_in4_3 = {io_validin64_51,io_in64_51}; // @[Cat.scala 30:58]
  assign ingress1_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 58:35]
  assign ingress1_13_clock = clock;
  assign ingress1_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign ingress1_13_io_in4_1 = {io_validin64_53,io_in64_53}; // @[Cat.scala 30:58]
  assign ingress1_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign ingress1_13_io_in4_3 = {io_validin64_55,io_in64_55}; // @[Cat.scala 30:58]
  assign ingress1_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 58:35]
  assign ingress1_14_clock = clock;
  assign ingress1_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign ingress1_14_io_in4_1 = {io_validin64_57,io_in64_57}; // @[Cat.scala 30:58]
  assign ingress1_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign ingress1_14_io_in4_3 = {io_validin64_59,io_in64_59}; // @[Cat.scala 30:58]
  assign ingress1_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 58:35]
  assign ingress1_15_clock = clock;
  assign ingress1_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign ingress1_15_io_in4_1 = {io_validin64_61,io_in64_61}; // @[Cat.scala 30:58]
  assign ingress1_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign ingress1_15_io_in4_3 = {io_validin64_63,io_in64_63}; // @[Cat.scala 30:58]
  assign ingress1_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 58:35]
  always @(posedge clock) begin
    addr <= io_addrin; // @[BuildingBlock.scala 42:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOSingress2(
  input          clock,
  input  [3:0]   io_in64_0,
  input  [3:0]   io_in64_1,
  input  [3:0]   io_in64_2,
  input  [3:0]   io_in64_3,
  input  [3:0]   io_in64_4,
  input  [3:0]   io_in64_5,
  input  [3:0]   io_in64_6,
  input  [3:0]   io_in64_7,
  input  [3:0]   io_in64_8,
  input  [3:0]   io_in64_9,
  input  [3:0]   io_in64_10,
  input  [3:0]   io_in64_11,
  input  [3:0]   io_in64_12,
  input  [3:0]   io_in64_13,
  input  [3:0]   io_in64_14,
  input  [3:0]   io_in64_15,
  input  [3:0]   io_in64_16,
  input  [3:0]   io_in64_17,
  input  [3:0]   io_in64_18,
  input  [3:0]   io_in64_19,
  input  [3:0]   io_in64_20,
  input  [3:0]   io_in64_21,
  input  [3:0]   io_in64_22,
  input  [3:0]   io_in64_23,
  input  [3:0]   io_in64_24,
  input  [3:0]   io_in64_25,
  input  [3:0]   io_in64_26,
  input  [3:0]   io_in64_27,
  input  [3:0]   io_in64_28,
  input  [3:0]   io_in64_29,
  input  [3:0]   io_in64_30,
  input  [3:0]   io_in64_31,
  input  [3:0]   io_in64_32,
  input  [3:0]   io_in64_33,
  input  [3:0]   io_in64_34,
  input  [3:0]   io_in64_35,
  input  [3:0]   io_in64_36,
  input  [3:0]   io_in64_37,
  input  [3:0]   io_in64_38,
  input  [3:0]   io_in64_39,
  input  [3:0]   io_in64_40,
  input  [3:0]   io_in64_41,
  input  [3:0]   io_in64_42,
  input  [3:0]   io_in64_43,
  input  [3:0]   io_in64_44,
  input  [3:0]   io_in64_45,
  input  [3:0]   io_in64_46,
  input  [3:0]   io_in64_47,
  input  [3:0]   io_in64_48,
  input  [3:0]   io_in64_49,
  input  [3:0]   io_in64_50,
  input  [3:0]   io_in64_51,
  input  [3:0]   io_in64_52,
  input  [3:0]   io_in64_53,
  input  [3:0]   io_in64_54,
  input  [3:0]   io_in64_55,
  input  [3:0]   io_in64_56,
  input  [3:0]   io_in64_57,
  input  [3:0]   io_in64_58,
  input  [3:0]   io_in64_59,
  input  [3:0]   io_in64_60,
  input  [3:0]   io_in64_61,
  input  [3:0]   io_in64_62,
  input  [3:0]   io_in64_63,
  input          io_validin64_0,
  input          io_validin64_1,
  input          io_validin64_2,
  input          io_validin64_3,
  input          io_validin64_4,
  input          io_validin64_5,
  input          io_validin64_6,
  input          io_validin64_7,
  input          io_validin64_8,
  input          io_validin64_9,
  input          io_validin64_10,
  input          io_validin64_11,
  input          io_validin64_12,
  input          io_validin64_13,
  input          io_validin64_14,
  input          io_validin64_15,
  input          io_validin64_16,
  input          io_validin64_17,
  input          io_validin64_18,
  input          io_validin64_19,
  input          io_validin64_20,
  input          io_validin64_21,
  input          io_validin64_22,
  input          io_validin64_23,
  input          io_validin64_24,
  input          io_validin64_25,
  input          io_validin64_26,
  input          io_validin64_27,
  input          io_validin64_28,
  input          io_validin64_29,
  input          io_validin64_30,
  input          io_validin64_31,
  input          io_validin64_32,
  input          io_validin64_33,
  input          io_validin64_34,
  input          io_validin64_35,
  input          io_validin64_36,
  input          io_validin64_37,
  input          io_validin64_38,
  input          io_validin64_39,
  input          io_validin64_40,
  input          io_validin64_41,
  input          io_validin64_42,
  input          io_validin64_43,
  input          io_validin64_44,
  input          io_validin64_45,
  input          io_validin64_46,
  input          io_validin64_47,
  input          io_validin64_48,
  input          io_validin64_49,
  input          io_validin64_50,
  input          io_validin64_51,
  input          io_validin64_52,
  input          io_validin64_53,
  input          io_validin64_54,
  input          io_validin64_55,
  input          io_validin64_56,
  input          io_validin64_57,
  input          io_validin64_58,
  input          io_validin64_59,
  input          io_validin64_60,
  input          io_validin64_61,
  input          io_validin64_62,
  input          io_validin64_63,
  input  [7:0]   io_addrin,
  output [3:0]   io_out64_0,
  output [3:0]   io_out64_1,
  output [3:0]   io_out64_2,
  output [3:0]   io_out64_3,
  output [3:0]   io_out64_4,
  output [3:0]   io_out64_5,
  output [3:0]   io_out64_6,
  output [3:0]   io_out64_7,
  output [3:0]   io_out64_8,
  output [3:0]   io_out64_9,
  output [3:0]   io_out64_10,
  output [3:0]   io_out64_11,
  output [3:0]   io_out64_12,
  output [3:0]   io_out64_13,
  output [3:0]   io_out64_14,
  output [3:0]   io_out64_15,
  output [3:0]   io_out64_16,
  output [3:0]   io_out64_17,
  output [3:0]   io_out64_18,
  output [3:0]   io_out64_19,
  output [3:0]   io_out64_20,
  output [3:0]   io_out64_21,
  output [3:0]   io_out64_22,
  output [3:0]   io_out64_23,
  output [3:0]   io_out64_24,
  output [3:0]   io_out64_25,
  output [3:0]   io_out64_26,
  output [3:0]   io_out64_27,
  output [3:0]   io_out64_28,
  output [3:0]   io_out64_29,
  output [3:0]   io_out64_30,
  output [3:0]   io_out64_31,
  output [3:0]   io_out64_32,
  output [3:0]   io_out64_33,
  output [3:0]   io_out64_34,
  output [3:0]   io_out64_35,
  output [3:0]   io_out64_36,
  output [3:0]   io_out64_37,
  output [3:0]   io_out64_38,
  output [3:0]   io_out64_39,
  output [3:0]   io_out64_40,
  output [3:0]   io_out64_41,
  output [3:0]   io_out64_42,
  output [3:0]   io_out64_43,
  output [3:0]   io_out64_44,
  output [3:0]   io_out64_45,
  output [3:0]   io_out64_46,
  output [3:0]   io_out64_47,
  output [3:0]   io_out64_48,
  output [3:0]   io_out64_49,
  output [3:0]   io_out64_50,
  output [3:0]   io_out64_51,
  output [3:0]   io_out64_52,
  output [3:0]   io_out64_53,
  output [3:0]   io_out64_54,
  output [3:0]   io_out64_55,
  output [3:0]   io_out64_56,
  output [3:0]   io_out64_57,
  output [3:0]   io_out64_58,
  output [3:0]   io_out64_59,
  output [3:0]   io_out64_60,
  output [3:0]   io_out64_61,
  output [3:0]   io_out64_62,
  output [3:0]   io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  ingress2_0_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_0_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_0_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_1_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_1_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_1_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_2_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_2_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_2_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_3_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_3_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_3_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_4_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_4_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_4_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_5_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_5_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_5_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_6_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_6_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_6_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_7_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_7_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_7_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_8_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_8_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_8_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_9_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_9_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_9_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_10_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_10_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_10_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_11_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_11_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_11_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_12_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_12_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_12_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_13_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_13_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_13_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_14_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_14_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_14_io_ctrl; // @[BuildingBlock.scala 74:52]
  wire  ingress2_15_clock; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_in4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_in4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_in4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_in4_3; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_out4_0; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_out4_1; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_out4_2; // @[BuildingBlock.scala 74:52]
  wire [4:0] ingress2_15_io_out4_3; // @[BuildingBlock.scala 74:52]
  wire [7:0] ingress2_15_io_ctrl; // @[BuildingBlock.scala 74:52]
  reg [7:0] addr; // @[BuildingBlock.scala 77:21]
  CLOScell4 ingress2_0 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_0_clock),
    .io_in4_0(ingress2_0_io_in4_0),
    .io_in4_1(ingress2_0_io_in4_1),
    .io_in4_2(ingress2_0_io_in4_2),
    .io_in4_3(ingress2_0_io_in4_3),
    .io_out4_0(ingress2_0_io_out4_0),
    .io_out4_1(ingress2_0_io_out4_1),
    .io_out4_2(ingress2_0_io_out4_2),
    .io_out4_3(ingress2_0_io_out4_3),
    .io_ctrl(ingress2_0_io_ctrl)
  );
  CLOScell4 ingress2_1 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_1_clock),
    .io_in4_0(ingress2_1_io_in4_0),
    .io_in4_1(ingress2_1_io_in4_1),
    .io_in4_2(ingress2_1_io_in4_2),
    .io_in4_3(ingress2_1_io_in4_3),
    .io_out4_0(ingress2_1_io_out4_0),
    .io_out4_1(ingress2_1_io_out4_1),
    .io_out4_2(ingress2_1_io_out4_2),
    .io_out4_3(ingress2_1_io_out4_3),
    .io_ctrl(ingress2_1_io_ctrl)
  );
  CLOScell4 ingress2_2 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_2_clock),
    .io_in4_0(ingress2_2_io_in4_0),
    .io_in4_1(ingress2_2_io_in4_1),
    .io_in4_2(ingress2_2_io_in4_2),
    .io_in4_3(ingress2_2_io_in4_3),
    .io_out4_0(ingress2_2_io_out4_0),
    .io_out4_1(ingress2_2_io_out4_1),
    .io_out4_2(ingress2_2_io_out4_2),
    .io_out4_3(ingress2_2_io_out4_3),
    .io_ctrl(ingress2_2_io_ctrl)
  );
  CLOScell4 ingress2_3 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_3_clock),
    .io_in4_0(ingress2_3_io_in4_0),
    .io_in4_1(ingress2_3_io_in4_1),
    .io_in4_2(ingress2_3_io_in4_2),
    .io_in4_3(ingress2_3_io_in4_3),
    .io_out4_0(ingress2_3_io_out4_0),
    .io_out4_1(ingress2_3_io_out4_1),
    .io_out4_2(ingress2_3_io_out4_2),
    .io_out4_3(ingress2_3_io_out4_3),
    .io_ctrl(ingress2_3_io_ctrl)
  );
  CLOScell4 ingress2_4 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_4_clock),
    .io_in4_0(ingress2_4_io_in4_0),
    .io_in4_1(ingress2_4_io_in4_1),
    .io_in4_2(ingress2_4_io_in4_2),
    .io_in4_3(ingress2_4_io_in4_3),
    .io_out4_0(ingress2_4_io_out4_0),
    .io_out4_1(ingress2_4_io_out4_1),
    .io_out4_2(ingress2_4_io_out4_2),
    .io_out4_3(ingress2_4_io_out4_3),
    .io_ctrl(ingress2_4_io_ctrl)
  );
  CLOScell4 ingress2_5 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_5_clock),
    .io_in4_0(ingress2_5_io_in4_0),
    .io_in4_1(ingress2_5_io_in4_1),
    .io_in4_2(ingress2_5_io_in4_2),
    .io_in4_3(ingress2_5_io_in4_3),
    .io_out4_0(ingress2_5_io_out4_0),
    .io_out4_1(ingress2_5_io_out4_1),
    .io_out4_2(ingress2_5_io_out4_2),
    .io_out4_3(ingress2_5_io_out4_3),
    .io_ctrl(ingress2_5_io_ctrl)
  );
  CLOScell4 ingress2_6 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_6_clock),
    .io_in4_0(ingress2_6_io_in4_0),
    .io_in4_1(ingress2_6_io_in4_1),
    .io_in4_2(ingress2_6_io_in4_2),
    .io_in4_3(ingress2_6_io_in4_3),
    .io_out4_0(ingress2_6_io_out4_0),
    .io_out4_1(ingress2_6_io_out4_1),
    .io_out4_2(ingress2_6_io_out4_2),
    .io_out4_3(ingress2_6_io_out4_3),
    .io_ctrl(ingress2_6_io_ctrl)
  );
  CLOScell4 ingress2_7 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_7_clock),
    .io_in4_0(ingress2_7_io_in4_0),
    .io_in4_1(ingress2_7_io_in4_1),
    .io_in4_2(ingress2_7_io_in4_2),
    .io_in4_3(ingress2_7_io_in4_3),
    .io_out4_0(ingress2_7_io_out4_0),
    .io_out4_1(ingress2_7_io_out4_1),
    .io_out4_2(ingress2_7_io_out4_2),
    .io_out4_3(ingress2_7_io_out4_3),
    .io_ctrl(ingress2_7_io_ctrl)
  );
  CLOScell4 ingress2_8 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_8_clock),
    .io_in4_0(ingress2_8_io_in4_0),
    .io_in4_1(ingress2_8_io_in4_1),
    .io_in4_2(ingress2_8_io_in4_2),
    .io_in4_3(ingress2_8_io_in4_3),
    .io_out4_0(ingress2_8_io_out4_0),
    .io_out4_1(ingress2_8_io_out4_1),
    .io_out4_2(ingress2_8_io_out4_2),
    .io_out4_3(ingress2_8_io_out4_3),
    .io_ctrl(ingress2_8_io_ctrl)
  );
  CLOScell4 ingress2_9 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_9_clock),
    .io_in4_0(ingress2_9_io_in4_0),
    .io_in4_1(ingress2_9_io_in4_1),
    .io_in4_2(ingress2_9_io_in4_2),
    .io_in4_3(ingress2_9_io_in4_3),
    .io_out4_0(ingress2_9_io_out4_0),
    .io_out4_1(ingress2_9_io_out4_1),
    .io_out4_2(ingress2_9_io_out4_2),
    .io_out4_3(ingress2_9_io_out4_3),
    .io_ctrl(ingress2_9_io_ctrl)
  );
  CLOScell4 ingress2_10 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_10_clock),
    .io_in4_0(ingress2_10_io_in4_0),
    .io_in4_1(ingress2_10_io_in4_1),
    .io_in4_2(ingress2_10_io_in4_2),
    .io_in4_3(ingress2_10_io_in4_3),
    .io_out4_0(ingress2_10_io_out4_0),
    .io_out4_1(ingress2_10_io_out4_1),
    .io_out4_2(ingress2_10_io_out4_2),
    .io_out4_3(ingress2_10_io_out4_3),
    .io_ctrl(ingress2_10_io_ctrl)
  );
  CLOScell4 ingress2_11 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_11_clock),
    .io_in4_0(ingress2_11_io_in4_0),
    .io_in4_1(ingress2_11_io_in4_1),
    .io_in4_2(ingress2_11_io_in4_2),
    .io_in4_3(ingress2_11_io_in4_3),
    .io_out4_0(ingress2_11_io_out4_0),
    .io_out4_1(ingress2_11_io_out4_1),
    .io_out4_2(ingress2_11_io_out4_2),
    .io_out4_3(ingress2_11_io_out4_3),
    .io_ctrl(ingress2_11_io_ctrl)
  );
  CLOScell4 ingress2_12 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_12_clock),
    .io_in4_0(ingress2_12_io_in4_0),
    .io_in4_1(ingress2_12_io_in4_1),
    .io_in4_2(ingress2_12_io_in4_2),
    .io_in4_3(ingress2_12_io_in4_3),
    .io_out4_0(ingress2_12_io_out4_0),
    .io_out4_1(ingress2_12_io_out4_1),
    .io_out4_2(ingress2_12_io_out4_2),
    .io_out4_3(ingress2_12_io_out4_3),
    .io_ctrl(ingress2_12_io_ctrl)
  );
  CLOScell4 ingress2_13 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_13_clock),
    .io_in4_0(ingress2_13_io_in4_0),
    .io_in4_1(ingress2_13_io_in4_1),
    .io_in4_2(ingress2_13_io_in4_2),
    .io_in4_3(ingress2_13_io_in4_3),
    .io_out4_0(ingress2_13_io_out4_0),
    .io_out4_1(ingress2_13_io_out4_1),
    .io_out4_2(ingress2_13_io_out4_2),
    .io_out4_3(ingress2_13_io_out4_3),
    .io_ctrl(ingress2_13_io_ctrl)
  );
  CLOScell4 ingress2_14 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_14_clock),
    .io_in4_0(ingress2_14_io_in4_0),
    .io_in4_1(ingress2_14_io_in4_1),
    .io_in4_2(ingress2_14_io_in4_2),
    .io_in4_3(ingress2_14_io_in4_3),
    .io_out4_0(ingress2_14_io_out4_0),
    .io_out4_1(ingress2_14_io_out4_1),
    .io_out4_2(ingress2_14_io_out4_2),
    .io_out4_3(ingress2_14_io_out4_3),
    .io_ctrl(ingress2_14_io_ctrl)
  );
  CLOScell4 ingress2_15 ( // @[BuildingBlock.scala 74:52]
    .clock(ingress2_15_clock),
    .io_in4_0(ingress2_15_io_in4_0),
    .io_in4_1(ingress2_15_io_in4_1),
    .io_in4_2(ingress2_15_io_in4_2),
    .io_in4_3(ingress2_15_io_in4_3),
    .io_out4_0(ingress2_15_io_out4_0),
    .io_out4_1(ingress2_15_io_out4_1),
    .io_out4_2(ingress2_15_io_out4_2),
    .io_out4_3(ingress2_15_io_out4_3),
    .io_ctrl(ingress2_15_io_ctrl)
  );
  assign io_out64_0 = ingress2_0_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_1 = ingress2_1_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_2 = ingress2_2_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_3 = ingress2_3_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_4 = ingress2_0_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_5 = ingress2_1_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_6 = ingress2_2_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_7 = ingress2_3_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_8 = ingress2_0_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_9 = ingress2_1_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_10 = ingress2_2_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_11 = ingress2_3_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_12 = ingress2_0_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_13 = ingress2_1_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_14 = ingress2_2_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_15 = ingress2_3_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_16 = ingress2_4_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_17 = ingress2_5_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_18 = ingress2_6_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_19 = ingress2_7_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_20 = ingress2_4_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_21 = ingress2_5_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_22 = ingress2_6_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_23 = ingress2_7_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_24 = ingress2_4_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_25 = ingress2_5_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_26 = ingress2_6_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_27 = ingress2_7_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_28 = ingress2_4_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_29 = ingress2_5_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_30 = ingress2_6_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_31 = ingress2_7_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_32 = ingress2_8_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_33 = ingress2_9_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_34 = ingress2_10_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_35 = ingress2_11_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_36 = ingress2_8_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_37 = ingress2_9_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_38 = ingress2_10_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_39 = ingress2_11_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_40 = ingress2_8_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_41 = ingress2_9_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_42 = ingress2_10_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_43 = ingress2_11_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_44 = ingress2_8_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_45 = ingress2_9_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_46 = ingress2_10_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_47 = ingress2_11_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_48 = ingress2_12_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_49 = ingress2_13_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_50 = ingress2_14_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_51 = ingress2_15_io_out4_0[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_52 = ingress2_12_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_53 = ingress2_13_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_54 = ingress2_14_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_55 = ingress2_15_io_out4_1[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_56 = ingress2_12_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_57 = ingress2_13_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_58 = ingress2_14_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_59 = ingress2_15_io_out4_2[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_60 = ingress2_12_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_61 = ingress2_13_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_62 = ingress2_14_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_out64_63 = ingress2_15_io_out4_3[3:0]; // @[BuildingBlock.scala 89:59]
  assign io_validout64_0 = ingress2_0_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_1 = ingress2_1_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_2 = ingress2_2_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_3 = ingress2_3_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_4 = ingress2_0_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_5 = ingress2_1_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_6 = ingress2_2_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_7 = ingress2_3_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_8 = ingress2_0_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_9 = ingress2_1_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_10 = ingress2_2_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_11 = ingress2_3_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_12 = ingress2_0_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_13 = ingress2_1_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_14 = ingress2_2_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_15 = ingress2_3_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_16 = ingress2_4_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_17 = ingress2_5_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_18 = ingress2_6_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_19 = ingress2_7_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_20 = ingress2_4_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_21 = ingress2_5_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_22 = ingress2_6_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_23 = ingress2_7_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_24 = ingress2_4_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_25 = ingress2_5_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_26 = ingress2_6_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_27 = ingress2_7_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_28 = ingress2_4_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_29 = ingress2_5_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_30 = ingress2_6_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_31 = ingress2_7_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_32 = ingress2_8_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_33 = ingress2_9_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_34 = ingress2_10_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_35 = ingress2_11_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_36 = ingress2_8_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_37 = ingress2_9_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_38 = ingress2_10_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_39 = ingress2_11_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_40 = ingress2_8_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_41 = ingress2_9_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_42 = ingress2_10_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_43 = ingress2_11_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_44 = ingress2_8_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_45 = ingress2_9_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_46 = ingress2_10_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_47 = ingress2_11_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_48 = ingress2_12_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_49 = ingress2_13_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_50 = ingress2_14_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_51 = ingress2_15_io_out4_0[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_52 = ingress2_12_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_53 = ingress2_13_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_54 = ingress2_14_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_55 = ingress2_15_io_out4_1[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_56 = ingress2_12_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_57 = ingress2_13_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_58 = ingress2_14_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_59 = ingress2_15_io_out4_2[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_60 = ingress2_12_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_61 = ingress2_13_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_62 = ingress2_14_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_validout64_63 = ingress2_15_io_out4_3[4]; // @[BuildingBlock.scala 90:64]
  assign io_addrout = addr; // @[BuildingBlock.scala 78:14]
  assign ingress2_0_clock = clock;
  assign ingress2_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign ingress2_0_io_in4_1 = {io_validin64_1,io_in64_1}; // @[Cat.scala 30:58]
  assign ingress2_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign ingress2_0_io_in4_3 = {io_validin64_3,io_in64_3}; // @[Cat.scala 30:58]
  assign ingress2_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 94:35]
  assign ingress2_1_clock = clock;
  assign ingress2_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign ingress2_1_io_in4_1 = {io_validin64_5,io_in64_5}; // @[Cat.scala 30:58]
  assign ingress2_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign ingress2_1_io_in4_3 = {io_validin64_7,io_in64_7}; // @[Cat.scala 30:58]
  assign ingress2_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 94:35]
  assign ingress2_2_clock = clock;
  assign ingress2_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign ingress2_2_io_in4_1 = {io_validin64_9,io_in64_9}; // @[Cat.scala 30:58]
  assign ingress2_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign ingress2_2_io_in4_3 = {io_validin64_11,io_in64_11}; // @[Cat.scala 30:58]
  assign ingress2_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 94:35]
  assign ingress2_3_clock = clock;
  assign ingress2_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign ingress2_3_io_in4_1 = {io_validin64_13,io_in64_13}; // @[Cat.scala 30:58]
  assign ingress2_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign ingress2_3_io_in4_3 = {io_validin64_15,io_in64_15}; // @[Cat.scala 30:58]
  assign ingress2_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 94:35]
  assign ingress2_4_clock = clock;
  assign ingress2_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign ingress2_4_io_in4_1 = {io_validin64_17,io_in64_17}; // @[Cat.scala 30:58]
  assign ingress2_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign ingress2_4_io_in4_3 = {io_validin64_19,io_in64_19}; // @[Cat.scala 30:58]
  assign ingress2_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 94:35]
  assign ingress2_5_clock = clock;
  assign ingress2_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign ingress2_5_io_in4_1 = {io_validin64_21,io_in64_21}; // @[Cat.scala 30:58]
  assign ingress2_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign ingress2_5_io_in4_3 = {io_validin64_23,io_in64_23}; // @[Cat.scala 30:58]
  assign ingress2_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 94:35]
  assign ingress2_6_clock = clock;
  assign ingress2_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign ingress2_6_io_in4_1 = {io_validin64_25,io_in64_25}; // @[Cat.scala 30:58]
  assign ingress2_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign ingress2_6_io_in4_3 = {io_validin64_27,io_in64_27}; // @[Cat.scala 30:58]
  assign ingress2_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 94:35]
  assign ingress2_7_clock = clock;
  assign ingress2_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign ingress2_7_io_in4_1 = {io_validin64_29,io_in64_29}; // @[Cat.scala 30:58]
  assign ingress2_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign ingress2_7_io_in4_3 = {io_validin64_31,io_in64_31}; // @[Cat.scala 30:58]
  assign ingress2_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 94:35]
  assign ingress2_8_clock = clock;
  assign ingress2_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign ingress2_8_io_in4_1 = {io_validin64_33,io_in64_33}; // @[Cat.scala 30:58]
  assign ingress2_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign ingress2_8_io_in4_3 = {io_validin64_35,io_in64_35}; // @[Cat.scala 30:58]
  assign ingress2_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 94:35]
  assign ingress2_9_clock = clock;
  assign ingress2_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign ingress2_9_io_in4_1 = {io_validin64_37,io_in64_37}; // @[Cat.scala 30:58]
  assign ingress2_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign ingress2_9_io_in4_3 = {io_validin64_39,io_in64_39}; // @[Cat.scala 30:58]
  assign ingress2_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 94:35]
  assign ingress2_10_clock = clock;
  assign ingress2_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign ingress2_10_io_in4_1 = {io_validin64_41,io_in64_41}; // @[Cat.scala 30:58]
  assign ingress2_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign ingress2_10_io_in4_3 = {io_validin64_43,io_in64_43}; // @[Cat.scala 30:58]
  assign ingress2_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 94:35]
  assign ingress2_11_clock = clock;
  assign ingress2_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign ingress2_11_io_in4_1 = {io_validin64_45,io_in64_45}; // @[Cat.scala 30:58]
  assign ingress2_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign ingress2_11_io_in4_3 = {io_validin64_47,io_in64_47}; // @[Cat.scala 30:58]
  assign ingress2_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 94:35]
  assign ingress2_12_clock = clock;
  assign ingress2_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign ingress2_12_io_in4_1 = {io_validin64_49,io_in64_49}; // @[Cat.scala 30:58]
  assign ingress2_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign ingress2_12_io_in4_3 = {io_validin64_51,io_in64_51}; // @[Cat.scala 30:58]
  assign ingress2_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 94:35]
  assign ingress2_13_clock = clock;
  assign ingress2_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign ingress2_13_io_in4_1 = {io_validin64_53,io_in64_53}; // @[Cat.scala 30:58]
  assign ingress2_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign ingress2_13_io_in4_3 = {io_validin64_55,io_in64_55}; // @[Cat.scala 30:58]
  assign ingress2_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 94:35]
  assign ingress2_14_clock = clock;
  assign ingress2_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign ingress2_14_io_in4_1 = {io_validin64_57,io_in64_57}; // @[Cat.scala 30:58]
  assign ingress2_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign ingress2_14_io_in4_3 = {io_validin64_59,io_in64_59}; // @[Cat.scala 30:58]
  assign ingress2_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 94:35]
  assign ingress2_15_clock = clock;
  assign ingress2_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign ingress2_15_io_in4_1 = {io_validin64_61,io_in64_61}; // @[Cat.scala 30:58]
  assign ingress2_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign ingress2_15_io_in4_3 = {io_validin64_63,io_in64_63}; // @[Cat.scala 30:58]
  assign ingress2_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 94:35]
  always @(posedge clock) begin
    addr <= io_addrin; // @[BuildingBlock.scala 77:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOSegress1(
  input          clock,
  input  [3:0]   io_in64_0,
  input  [3:0]   io_in64_1,
  input  [3:0]   io_in64_2,
  input  [3:0]   io_in64_3,
  input  [3:0]   io_in64_4,
  input  [3:0]   io_in64_5,
  input  [3:0]   io_in64_6,
  input  [3:0]   io_in64_7,
  input  [3:0]   io_in64_8,
  input  [3:0]   io_in64_9,
  input  [3:0]   io_in64_10,
  input  [3:0]   io_in64_11,
  input  [3:0]   io_in64_12,
  input  [3:0]   io_in64_13,
  input  [3:0]   io_in64_14,
  input  [3:0]   io_in64_15,
  input  [3:0]   io_in64_16,
  input  [3:0]   io_in64_17,
  input  [3:0]   io_in64_18,
  input  [3:0]   io_in64_19,
  input  [3:0]   io_in64_20,
  input  [3:0]   io_in64_21,
  input  [3:0]   io_in64_22,
  input  [3:0]   io_in64_23,
  input  [3:0]   io_in64_24,
  input  [3:0]   io_in64_25,
  input  [3:0]   io_in64_26,
  input  [3:0]   io_in64_27,
  input  [3:0]   io_in64_28,
  input  [3:0]   io_in64_29,
  input  [3:0]   io_in64_30,
  input  [3:0]   io_in64_31,
  input  [3:0]   io_in64_32,
  input  [3:0]   io_in64_33,
  input  [3:0]   io_in64_34,
  input  [3:0]   io_in64_35,
  input  [3:0]   io_in64_36,
  input  [3:0]   io_in64_37,
  input  [3:0]   io_in64_38,
  input  [3:0]   io_in64_39,
  input  [3:0]   io_in64_40,
  input  [3:0]   io_in64_41,
  input  [3:0]   io_in64_42,
  input  [3:0]   io_in64_43,
  input  [3:0]   io_in64_44,
  input  [3:0]   io_in64_45,
  input  [3:0]   io_in64_46,
  input  [3:0]   io_in64_47,
  input  [3:0]   io_in64_48,
  input  [3:0]   io_in64_49,
  input  [3:0]   io_in64_50,
  input  [3:0]   io_in64_51,
  input  [3:0]   io_in64_52,
  input  [3:0]   io_in64_53,
  input  [3:0]   io_in64_54,
  input  [3:0]   io_in64_55,
  input  [3:0]   io_in64_56,
  input  [3:0]   io_in64_57,
  input  [3:0]   io_in64_58,
  input  [3:0]   io_in64_59,
  input  [3:0]   io_in64_60,
  input  [3:0]   io_in64_61,
  input  [3:0]   io_in64_62,
  input  [3:0]   io_in64_63,
  input          io_validin64_0,
  input          io_validin64_1,
  input          io_validin64_2,
  input          io_validin64_3,
  input          io_validin64_4,
  input          io_validin64_5,
  input          io_validin64_6,
  input          io_validin64_7,
  input          io_validin64_8,
  input          io_validin64_9,
  input          io_validin64_10,
  input          io_validin64_11,
  input          io_validin64_12,
  input          io_validin64_13,
  input          io_validin64_14,
  input          io_validin64_15,
  input          io_validin64_16,
  input          io_validin64_17,
  input          io_validin64_18,
  input          io_validin64_19,
  input          io_validin64_20,
  input          io_validin64_21,
  input          io_validin64_22,
  input          io_validin64_23,
  input          io_validin64_24,
  input          io_validin64_25,
  input          io_validin64_26,
  input          io_validin64_27,
  input          io_validin64_28,
  input          io_validin64_29,
  input          io_validin64_30,
  input          io_validin64_31,
  input          io_validin64_32,
  input          io_validin64_33,
  input          io_validin64_34,
  input          io_validin64_35,
  input          io_validin64_36,
  input          io_validin64_37,
  input          io_validin64_38,
  input          io_validin64_39,
  input          io_validin64_40,
  input          io_validin64_41,
  input          io_validin64_42,
  input          io_validin64_43,
  input          io_validin64_44,
  input          io_validin64_45,
  input          io_validin64_46,
  input          io_validin64_47,
  input          io_validin64_48,
  input          io_validin64_49,
  input          io_validin64_50,
  input          io_validin64_51,
  input          io_validin64_52,
  input          io_validin64_53,
  input          io_validin64_54,
  input          io_validin64_55,
  input          io_validin64_56,
  input          io_validin64_57,
  input          io_validin64_58,
  input          io_validin64_59,
  input          io_validin64_60,
  input          io_validin64_61,
  input          io_validin64_62,
  input          io_validin64_63,
  input  [7:0]   io_addrin,
  output [3:0]   io_out64_0,
  output [3:0]   io_out64_1,
  output [3:0]   io_out64_2,
  output [3:0]   io_out64_3,
  output [3:0]   io_out64_4,
  output [3:0]   io_out64_5,
  output [3:0]   io_out64_6,
  output [3:0]   io_out64_7,
  output [3:0]   io_out64_8,
  output [3:0]   io_out64_9,
  output [3:0]   io_out64_10,
  output [3:0]   io_out64_11,
  output [3:0]   io_out64_12,
  output [3:0]   io_out64_13,
  output [3:0]   io_out64_14,
  output [3:0]   io_out64_15,
  output [3:0]   io_out64_16,
  output [3:0]   io_out64_17,
  output [3:0]   io_out64_18,
  output [3:0]   io_out64_19,
  output [3:0]   io_out64_20,
  output [3:0]   io_out64_21,
  output [3:0]   io_out64_22,
  output [3:0]   io_out64_23,
  output [3:0]   io_out64_24,
  output [3:0]   io_out64_25,
  output [3:0]   io_out64_26,
  output [3:0]   io_out64_27,
  output [3:0]   io_out64_28,
  output [3:0]   io_out64_29,
  output [3:0]   io_out64_30,
  output [3:0]   io_out64_31,
  output [3:0]   io_out64_32,
  output [3:0]   io_out64_33,
  output [3:0]   io_out64_34,
  output [3:0]   io_out64_35,
  output [3:0]   io_out64_36,
  output [3:0]   io_out64_37,
  output [3:0]   io_out64_38,
  output [3:0]   io_out64_39,
  output [3:0]   io_out64_40,
  output [3:0]   io_out64_41,
  output [3:0]   io_out64_42,
  output [3:0]   io_out64_43,
  output [3:0]   io_out64_44,
  output [3:0]   io_out64_45,
  output [3:0]   io_out64_46,
  output [3:0]   io_out64_47,
  output [3:0]   io_out64_48,
  output [3:0]   io_out64_49,
  output [3:0]   io_out64_50,
  output [3:0]   io_out64_51,
  output [3:0]   io_out64_52,
  output [3:0]   io_out64_53,
  output [3:0]   io_out64_54,
  output [3:0]   io_out64_55,
  output [3:0]   io_out64_56,
  output [3:0]   io_out64_57,
  output [3:0]   io_out64_58,
  output [3:0]   io_out64_59,
  output [3:0]   io_out64_60,
  output [3:0]   io_out64_61,
  output [3:0]   io_out64_62,
  output [3:0]   io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  egress1_0_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_0_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_0_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_1_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_1_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_1_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_2_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_2_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_2_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_3_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_3_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_3_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_4_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_4_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_4_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_5_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_5_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_5_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_6_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_6_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_6_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_7_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_7_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_7_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_8_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_8_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_8_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_9_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_9_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_9_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_10_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_10_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_10_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_11_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_11_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_11_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_12_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_12_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_12_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_13_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_13_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_13_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_14_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_14_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_14_io_ctrl; // @[BuildingBlock.scala 147:51]
  wire  egress1_15_clock; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_in4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_in4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_in4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_in4_3; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_out4_0; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_out4_1; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_out4_2; // @[BuildingBlock.scala 147:51]
  wire [4:0] egress1_15_io_out4_3; // @[BuildingBlock.scala 147:51]
  wire [7:0] egress1_15_io_ctrl; // @[BuildingBlock.scala 147:51]
  reg [7:0] addr; // @[BuildingBlock.scala 150:21]
  CLOScell4 egress1_0 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_0_clock),
    .io_in4_0(egress1_0_io_in4_0),
    .io_in4_1(egress1_0_io_in4_1),
    .io_in4_2(egress1_0_io_in4_2),
    .io_in4_3(egress1_0_io_in4_3),
    .io_out4_0(egress1_0_io_out4_0),
    .io_out4_1(egress1_0_io_out4_1),
    .io_out4_2(egress1_0_io_out4_2),
    .io_out4_3(egress1_0_io_out4_3),
    .io_ctrl(egress1_0_io_ctrl)
  );
  CLOScell4 egress1_1 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_1_clock),
    .io_in4_0(egress1_1_io_in4_0),
    .io_in4_1(egress1_1_io_in4_1),
    .io_in4_2(egress1_1_io_in4_2),
    .io_in4_3(egress1_1_io_in4_3),
    .io_out4_0(egress1_1_io_out4_0),
    .io_out4_1(egress1_1_io_out4_1),
    .io_out4_2(egress1_1_io_out4_2),
    .io_out4_3(egress1_1_io_out4_3),
    .io_ctrl(egress1_1_io_ctrl)
  );
  CLOScell4 egress1_2 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_2_clock),
    .io_in4_0(egress1_2_io_in4_0),
    .io_in4_1(egress1_2_io_in4_1),
    .io_in4_2(egress1_2_io_in4_2),
    .io_in4_3(egress1_2_io_in4_3),
    .io_out4_0(egress1_2_io_out4_0),
    .io_out4_1(egress1_2_io_out4_1),
    .io_out4_2(egress1_2_io_out4_2),
    .io_out4_3(egress1_2_io_out4_3),
    .io_ctrl(egress1_2_io_ctrl)
  );
  CLOScell4 egress1_3 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_3_clock),
    .io_in4_0(egress1_3_io_in4_0),
    .io_in4_1(egress1_3_io_in4_1),
    .io_in4_2(egress1_3_io_in4_2),
    .io_in4_3(egress1_3_io_in4_3),
    .io_out4_0(egress1_3_io_out4_0),
    .io_out4_1(egress1_3_io_out4_1),
    .io_out4_2(egress1_3_io_out4_2),
    .io_out4_3(egress1_3_io_out4_3),
    .io_ctrl(egress1_3_io_ctrl)
  );
  CLOScell4 egress1_4 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_4_clock),
    .io_in4_0(egress1_4_io_in4_0),
    .io_in4_1(egress1_4_io_in4_1),
    .io_in4_2(egress1_4_io_in4_2),
    .io_in4_3(egress1_4_io_in4_3),
    .io_out4_0(egress1_4_io_out4_0),
    .io_out4_1(egress1_4_io_out4_1),
    .io_out4_2(egress1_4_io_out4_2),
    .io_out4_3(egress1_4_io_out4_3),
    .io_ctrl(egress1_4_io_ctrl)
  );
  CLOScell4 egress1_5 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_5_clock),
    .io_in4_0(egress1_5_io_in4_0),
    .io_in4_1(egress1_5_io_in4_1),
    .io_in4_2(egress1_5_io_in4_2),
    .io_in4_3(egress1_5_io_in4_3),
    .io_out4_0(egress1_5_io_out4_0),
    .io_out4_1(egress1_5_io_out4_1),
    .io_out4_2(egress1_5_io_out4_2),
    .io_out4_3(egress1_5_io_out4_3),
    .io_ctrl(egress1_5_io_ctrl)
  );
  CLOScell4 egress1_6 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_6_clock),
    .io_in4_0(egress1_6_io_in4_0),
    .io_in4_1(egress1_6_io_in4_1),
    .io_in4_2(egress1_6_io_in4_2),
    .io_in4_3(egress1_6_io_in4_3),
    .io_out4_0(egress1_6_io_out4_0),
    .io_out4_1(egress1_6_io_out4_1),
    .io_out4_2(egress1_6_io_out4_2),
    .io_out4_3(egress1_6_io_out4_3),
    .io_ctrl(egress1_6_io_ctrl)
  );
  CLOScell4 egress1_7 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_7_clock),
    .io_in4_0(egress1_7_io_in4_0),
    .io_in4_1(egress1_7_io_in4_1),
    .io_in4_2(egress1_7_io_in4_2),
    .io_in4_3(egress1_7_io_in4_3),
    .io_out4_0(egress1_7_io_out4_0),
    .io_out4_1(egress1_7_io_out4_1),
    .io_out4_2(egress1_7_io_out4_2),
    .io_out4_3(egress1_7_io_out4_3),
    .io_ctrl(egress1_7_io_ctrl)
  );
  CLOScell4 egress1_8 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_8_clock),
    .io_in4_0(egress1_8_io_in4_0),
    .io_in4_1(egress1_8_io_in4_1),
    .io_in4_2(egress1_8_io_in4_2),
    .io_in4_3(egress1_8_io_in4_3),
    .io_out4_0(egress1_8_io_out4_0),
    .io_out4_1(egress1_8_io_out4_1),
    .io_out4_2(egress1_8_io_out4_2),
    .io_out4_3(egress1_8_io_out4_3),
    .io_ctrl(egress1_8_io_ctrl)
  );
  CLOScell4 egress1_9 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_9_clock),
    .io_in4_0(egress1_9_io_in4_0),
    .io_in4_1(egress1_9_io_in4_1),
    .io_in4_2(egress1_9_io_in4_2),
    .io_in4_3(egress1_9_io_in4_3),
    .io_out4_0(egress1_9_io_out4_0),
    .io_out4_1(egress1_9_io_out4_1),
    .io_out4_2(egress1_9_io_out4_2),
    .io_out4_3(egress1_9_io_out4_3),
    .io_ctrl(egress1_9_io_ctrl)
  );
  CLOScell4 egress1_10 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_10_clock),
    .io_in4_0(egress1_10_io_in4_0),
    .io_in4_1(egress1_10_io_in4_1),
    .io_in4_2(egress1_10_io_in4_2),
    .io_in4_3(egress1_10_io_in4_3),
    .io_out4_0(egress1_10_io_out4_0),
    .io_out4_1(egress1_10_io_out4_1),
    .io_out4_2(egress1_10_io_out4_2),
    .io_out4_3(egress1_10_io_out4_3),
    .io_ctrl(egress1_10_io_ctrl)
  );
  CLOScell4 egress1_11 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_11_clock),
    .io_in4_0(egress1_11_io_in4_0),
    .io_in4_1(egress1_11_io_in4_1),
    .io_in4_2(egress1_11_io_in4_2),
    .io_in4_3(egress1_11_io_in4_3),
    .io_out4_0(egress1_11_io_out4_0),
    .io_out4_1(egress1_11_io_out4_1),
    .io_out4_2(egress1_11_io_out4_2),
    .io_out4_3(egress1_11_io_out4_3),
    .io_ctrl(egress1_11_io_ctrl)
  );
  CLOScell4 egress1_12 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_12_clock),
    .io_in4_0(egress1_12_io_in4_0),
    .io_in4_1(egress1_12_io_in4_1),
    .io_in4_2(egress1_12_io_in4_2),
    .io_in4_3(egress1_12_io_in4_3),
    .io_out4_0(egress1_12_io_out4_0),
    .io_out4_1(egress1_12_io_out4_1),
    .io_out4_2(egress1_12_io_out4_2),
    .io_out4_3(egress1_12_io_out4_3),
    .io_ctrl(egress1_12_io_ctrl)
  );
  CLOScell4 egress1_13 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_13_clock),
    .io_in4_0(egress1_13_io_in4_0),
    .io_in4_1(egress1_13_io_in4_1),
    .io_in4_2(egress1_13_io_in4_2),
    .io_in4_3(egress1_13_io_in4_3),
    .io_out4_0(egress1_13_io_out4_0),
    .io_out4_1(egress1_13_io_out4_1),
    .io_out4_2(egress1_13_io_out4_2),
    .io_out4_3(egress1_13_io_out4_3),
    .io_ctrl(egress1_13_io_ctrl)
  );
  CLOScell4 egress1_14 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_14_clock),
    .io_in4_0(egress1_14_io_in4_0),
    .io_in4_1(egress1_14_io_in4_1),
    .io_in4_2(egress1_14_io_in4_2),
    .io_in4_3(egress1_14_io_in4_3),
    .io_out4_0(egress1_14_io_out4_0),
    .io_out4_1(egress1_14_io_out4_1),
    .io_out4_2(egress1_14_io_out4_2),
    .io_out4_3(egress1_14_io_out4_3),
    .io_ctrl(egress1_14_io_ctrl)
  );
  CLOScell4 egress1_15 ( // @[BuildingBlock.scala 147:51]
    .clock(egress1_15_clock),
    .io_in4_0(egress1_15_io_in4_0),
    .io_in4_1(egress1_15_io_in4_1),
    .io_in4_2(egress1_15_io_in4_2),
    .io_in4_3(egress1_15_io_in4_3),
    .io_out4_0(egress1_15_io_out4_0),
    .io_out4_1(egress1_15_io_out4_1),
    .io_out4_2(egress1_15_io_out4_2),
    .io_out4_3(egress1_15_io_out4_3),
    .io_ctrl(egress1_15_io_ctrl)
  );
  assign io_out64_0 = egress1_0_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_1 = egress1_4_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_2 = egress1_8_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_3 = egress1_12_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_4 = egress1_0_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_5 = egress1_4_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_6 = egress1_8_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_7 = egress1_12_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_8 = egress1_0_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_9 = egress1_4_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_10 = egress1_8_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_11 = egress1_12_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_12 = egress1_0_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_13 = egress1_4_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_14 = egress1_8_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_15 = egress1_12_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_16 = egress1_1_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_17 = egress1_5_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_18 = egress1_9_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_19 = egress1_13_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_20 = egress1_1_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_21 = egress1_5_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_22 = egress1_9_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_23 = egress1_13_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_24 = egress1_1_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_25 = egress1_5_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_26 = egress1_9_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_27 = egress1_13_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_28 = egress1_1_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_29 = egress1_5_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_30 = egress1_9_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_31 = egress1_13_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_32 = egress1_2_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_33 = egress1_6_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_34 = egress1_10_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_35 = egress1_14_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_36 = egress1_2_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_37 = egress1_6_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_38 = egress1_10_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_39 = egress1_14_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_40 = egress1_2_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_41 = egress1_6_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_42 = egress1_10_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_43 = egress1_14_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_44 = egress1_2_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_45 = egress1_6_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_46 = egress1_10_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_47 = egress1_14_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_48 = egress1_3_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_49 = egress1_7_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_50 = egress1_11_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_51 = egress1_15_io_out4_0[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_52 = egress1_3_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_53 = egress1_7_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_54 = egress1_11_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_55 = egress1_15_io_out4_1[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_56 = egress1_3_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_57 = egress1_7_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_58 = egress1_11_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_59 = egress1_15_io_out4_2[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_60 = egress1_3_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_61 = egress1_7_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_62 = egress1_11_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_out64_63 = egress1_15_io_out4_3[3:0]; // @[BuildingBlock.scala 169:58]
  assign io_validout64_0 = egress1_0_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_1 = egress1_4_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_2 = egress1_8_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_3 = egress1_12_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_4 = egress1_0_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_5 = egress1_4_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_6 = egress1_8_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_7 = egress1_12_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_8 = egress1_0_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_9 = egress1_4_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_10 = egress1_8_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_11 = egress1_12_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_12 = egress1_0_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_13 = egress1_4_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_14 = egress1_8_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_15 = egress1_12_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_16 = egress1_1_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_17 = egress1_5_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_18 = egress1_9_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_19 = egress1_13_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_20 = egress1_1_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_21 = egress1_5_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_22 = egress1_9_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_23 = egress1_13_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_24 = egress1_1_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_25 = egress1_5_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_26 = egress1_9_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_27 = egress1_13_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_28 = egress1_1_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_29 = egress1_5_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_30 = egress1_9_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_31 = egress1_13_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_32 = egress1_2_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_33 = egress1_6_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_34 = egress1_10_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_35 = egress1_14_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_36 = egress1_2_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_37 = egress1_6_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_38 = egress1_10_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_39 = egress1_14_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_40 = egress1_2_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_41 = egress1_6_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_42 = egress1_10_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_43 = egress1_14_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_44 = egress1_2_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_45 = egress1_6_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_46 = egress1_10_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_47 = egress1_14_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_48 = egress1_3_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_49 = egress1_7_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_50 = egress1_11_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_51 = egress1_15_io_out4_0[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_52 = egress1_3_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_53 = egress1_7_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_54 = egress1_11_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_55 = egress1_15_io_out4_1[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_56 = egress1_3_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_57 = egress1_7_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_58 = egress1_11_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_59 = egress1_15_io_out4_2[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_60 = egress1_3_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_61 = egress1_7_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_62 = egress1_11_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_validout64_63 = egress1_15_io_out4_3[4]; // @[BuildingBlock.scala 170:63]
  assign io_addrout = addr; // @[BuildingBlock.scala 151:14]
  assign egress1_0_clock = clock;
  assign egress1_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign egress1_0_io_in4_1 = {io_validin64_1,io_in64_1}; // @[Cat.scala 30:58]
  assign egress1_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign egress1_0_io_in4_3 = {io_validin64_3,io_in64_3}; // @[Cat.scala 30:58]
  assign egress1_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 176:34]
  assign egress1_1_clock = clock;
  assign egress1_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign egress1_1_io_in4_1 = {io_validin64_5,io_in64_5}; // @[Cat.scala 30:58]
  assign egress1_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign egress1_1_io_in4_3 = {io_validin64_7,io_in64_7}; // @[Cat.scala 30:58]
  assign egress1_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 176:34]
  assign egress1_2_clock = clock;
  assign egress1_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign egress1_2_io_in4_1 = {io_validin64_9,io_in64_9}; // @[Cat.scala 30:58]
  assign egress1_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign egress1_2_io_in4_3 = {io_validin64_11,io_in64_11}; // @[Cat.scala 30:58]
  assign egress1_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 176:34]
  assign egress1_3_clock = clock;
  assign egress1_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign egress1_3_io_in4_1 = {io_validin64_13,io_in64_13}; // @[Cat.scala 30:58]
  assign egress1_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign egress1_3_io_in4_3 = {io_validin64_15,io_in64_15}; // @[Cat.scala 30:58]
  assign egress1_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 176:34]
  assign egress1_4_clock = clock;
  assign egress1_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign egress1_4_io_in4_1 = {io_validin64_17,io_in64_17}; // @[Cat.scala 30:58]
  assign egress1_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign egress1_4_io_in4_3 = {io_validin64_19,io_in64_19}; // @[Cat.scala 30:58]
  assign egress1_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 176:34]
  assign egress1_5_clock = clock;
  assign egress1_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign egress1_5_io_in4_1 = {io_validin64_21,io_in64_21}; // @[Cat.scala 30:58]
  assign egress1_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign egress1_5_io_in4_3 = {io_validin64_23,io_in64_23}; // @[Cat.scala 30:58]
  assign egress1_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 176:34]
  assign egress1_6_clock = clock;
  assign egress1_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign egress1_6_io_in4_1 = {io_validin64_25,io_in64_25}; // @[Cat.scala 30:58]
  assign egress1_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign egress1_6_io_in4_3 = {io_validin64_27,io_in64_27}; // @[Cat.scala 30:58]
  assign egress1_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 176:34]
  assign egress1_7_clock = clock;
  assign egress1_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign egress1_7_io_in4_1 = {io_validin64_29,io_in64_29}; // @[Cat.scala 30:58]
  assign egress1_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign egress1_7_io_in4_3 = {io_validin64_31,io_in64_31}; // @[Cat.scala 30:58]
  assign egress1_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 176:34]
  assign egress1_8_clock = clock;
  assign egress1_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign egress1_8_io_in4_1 = {io_validin64_33,io_in64_33}; // @[Cat.scala 30:58]
  assign egress1_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign egress1_8_io_in4_3 = {io_validin64_35,io_in64_35}; // @[Cat.scala 30:58]
  assign egress1_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 176:34]
  assign egress1_9_clock = clock;
  assign egress1_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign egress1_9_io_in4_1 = {io_validin64_37,io_in64_37}; // @[Cat.scala 30:58]
  assign egress1_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign egress1_9_io_in4_3 = {io_validin64_39,io_in64_39}; // @[Cat.scala 30:58]
  assign egress1_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 176:34]
  assign egress1_10_clock = clock;
  assign egress1_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign egress1_10_io_in4_1 = {io_validin64_41,io_in64_41}; // @[Cat.scala 30:58]
  assign egress1_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign egress1_10_io_in4_3 = {io_validin64_43,io_in64_43}; // @[Cat.scala 30:58]
  assign egress1_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 176:34]
  assign egress1_11_clock = clock;
  assign egress1_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign egress1_11_io_in4_1 = {io_validin64_45,io_in64_45}; // @[Cat.scala 30:58]
  assign egress1_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign egress1_11_io_in4_3 = {io_validin64_47,io_in64_47}; // @[Cat.scala 30:58]
  assign egress1_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 176:34]
  assign egress1_12_clock = clock;
  assign egress1_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign egress1_12_io_in4_1 = {io_validin64_49,io_in64_49}; // @[Cat.scala 30:58]
  assign egress1_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign egress1_12_io_in4_3 = {io_validin64_51,io_in64_51}; // @[Cat.scala 30:58]
  assign egress1_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 176:34]
  assign egress1_13_clock = clock;
  assign egress1_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign egress1_13_io_in4_1 = {io_validin64_53,io_in64_53}; // @[Cat.scala 30:58]
  assign egress1_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign egress1_13_io_in4_3 = {io_validin64_55,io_in64_55}; // @[Cat.scala 30:58]
  assign egress1_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 176:34]
  assign egress1_14_clock = clock;
  assign egress1_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign egress1_14_io_in4_1 = {io_validin64_57,io_in64_57}; // @[Cat.scala 30:58]
  assign egress1_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign egress1_14_io_in4_3 = {io_validin64_59,io_in64_59}; // @[Cat.scala 30:58]
  assign egress1_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 176:34]
  assign egress1_15_clock = clock;
  assign egress1_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign egress1_15_io_in4_1 = {io_validin64_61,io_in64_61}; // @[Cat.scala 30:58]
  assign egress1_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign egress1_15_io_in4_3 = {io_validin64_63,io_in64_63}; // @[Cat.scala 30:58]
  assign egress1_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 176:34]
  always @(posedge clock) begin
    addr <= io_addrin; // @[BuildingBlock.scala 150:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module CLOSegress2(
  input          clock,
  input  [3:0]   io_in64_0,
  input  [3:0]   io_in64_1,
  input  [3:0]   io_in64_2,
  input  [3:0]   io_in64_3,
  input  [3:0]   io_in64_4,
  input  [3:0]   io_in64_5,
  input  [3:0]   io_in64_6,
  input  [3:0]   io_in64_7,
  input  [3:0]   io_in64_8,
  input  [3:0]   io_in64_9,
  input  [3:0]   io_in64_10,
  input  [3:0]   io_in64_11,
  input  [3:0]   io_in64_12,
  input  [3:0]   io_in64_13,
  input  [3:0]   io_in64_14,
  input  [3:0]   io_in64_15,
  input  [3:0]   io_in64_16,
  input  [3:0]   io_in64_17,
  input  [3:0]   io_in64_18,
  input  [3:0]   io_in64_19,
  input  [3:0]   io_in64_20,
  input  [3:0]   io_in64_21,
  input  [3:0]   io_in64_22,
  input  [3:0]   io_in64_23,
  input  [3:0]   io_in64_24,
  input  [3:0]   io_in64_25,
  input  [3:0]   io_in64_26,
  input  [3:0]   io_in64_27,
  input  [3:0]   io_in64_28,
  input  [3:0]   io_in64_29,
  input  [3:0]   io_in64_30,
  input  [3:0]   io_in64_31,
  input  [3:0]   io_in64_32,
  input  [3:0]   io_in64_33,
  input  [3:0]   io_in64_34,
  input  [3:0]   io_in64_35,
  input  [3:0]   io_in64_36,
  input  [3:0]   io_in64_37,
  input  [3:0]   io_in64_38,
  input  [3:0]   io_in64_39,
  input  [3:0]   io_in64_40,
  input  [3:0]   io_in64_41,
  input  [3:0]   io_in64_42,
  input  [3:0]   io_in64_43,
  input  [3:0]   io_in64_44,
  input  [3:0]   io_in64_45,
  input  [3:0]   io_in64_46,
  input  [3:0]   io_in64_47,
  input  [3:0]   io_in64_48,
  input  [3:0]   io_in64_49,
  input  [3:0]   io_in64_50,
  input  [3:0]   io_in64_51,
  input  [3:0]   io_in64_52,
  input  [3:0]   io_in64_53,
  input  [3:0]   io_in64_54,
  input  [3:0]   io_in64_55,
  input  [3:0]   io_in64_56,
  input  [3:0]   io_in64_57,
  input  [3:0]   io_in64_58,
  input  [3:0]   io_in64_59,
  input  [3:0]   io_in64_60,
  input  [3:0]   io_in64_61,
  input  [3:0]   io_in64_62,
  input  [3:0]   io_in64_63,
  input          io_validin64_0,
  input          io_validin64_1,
  input          io_validin64_2,
  input          io_validin64_3,
  input          io_validin64_4,
  input          io_validin64_5,
  input          io_validin64_6,
  input          io_validin64_7,
  input          io_validin64_8,
  input          io_validin64_9,
  input          io_validin64_10,
  input          io_validin64_11,
  input          io_validin64_12,
  input          io_validin64_13,
  input          io_validin64_14,
  input          io_validin64_15,
  input          io_validin64_16,
  input          io_validin64_17,
  input          io_validin64_18,
  input          io_validin64_19,
  input          io_validin64_20,
  input          io_validin64_21,
  input          io_validin64_22,
  input          io_validin64_23,
  input          io_validin64_24,
  input          io_validin64_25,
  input          io_validin64_26,
  input          io_validin64_27,
  input          io_validin64_28,
  input          io_validin64_29,
  input          io_validin64_30,
  input          io_validin64_31,
  input          io_validin64_32,
  input          io_validin64_33,
  input          io_validin64_34,
  input          io_validin64_35,
  input          io_validin64_36,
  input          io_validin64_37,
  input          io_validin64_38,
  input          io_validin64_39,
  input          io_validin64_40,
  input          io_validin64_41,
  input          io_validin64_42,
  input          io_validin64_43,
  input          io_validin64_44,
  input          io_validin64_45,
  input          io_validin64_46,
  input          io_validin64_47,
  input          io_validin64_48,
  input          io_validin64_49,
  input          io_validin64_50,
  input          io_validin64_51,
  input          io_validin64_52,
  input          io_validin64_53,
  input          io_validin64_54,
  input          io_validin64_55,
  input          io_validin64_56,
  input          io_validin64_57,
  input          io_validin64_58,
  input          io_validin64_59,
  input          io_validin64_60,
  input          io_validin64_61,
  input          io_validin64_62,
  input          io_validin64_63,
  input  [7:0]   io_addrin,
  output [3:0]   io_out64_0,
  output [3:0]   io_out64_1,
  output [3:0]   io_out64_2,
  output [3:0]   io_out64_3,
  output [3:0]   io_out64_4,
  output [3:0]   io_out64_5,
  output [3:0]   io_out64_6,
  output [3:0]   io_out64_7,
  output [3:0]   io_out64_8,
  output [3:0]   io_out64_9,
  output [3:0]   io_out64_10,
  output [3:0]   io_out64_11,
  output [3:0]   io_out64_12,
  output [3:0]   io_out64_13,
  output [3:0]   io_out64_14,
  output [3:0]   io_out64_15,
  output [3:0]   io_out64_16,
  output [3:0]   io_out64_17,
  output [3:0]   io_out64_18,
  output [3:0]   io_out64_19,
  output [3:0]   io_out64_20,
  output [3:0]   io_out64_21,
  output [3:0]   io_out64_22,
  output [3:0]   io_out64_23,
  output [3:0]   io_out64_24,
  output [3:0]   io_out64_25,
  output [3:0]   io_out64_26,
  output [3:0]   io_out64_27,
  output [3:0]   io_out64_28,
  output [3:0]   io_out64_29,
  output [3:0]   io_out64_30,
  output [3:0]   io_out64_31,
  output [3:0]   io_out64_32,
  output [3:0]   io_out64_33,
  output [3:0]   io_out64_34,
  output [3:0]   io_out64_35,
  output [3:0]   io_out64_36,
  output [3:0]   io_out64_37,
  output [3:0]   io_out64_38,
  output [3:0]   io_out64_39,
  output [3:0]   io_out64_40,
  output [3:0]   io_out64_41,
  output [3:0]   io_out64_42,
  output [3:0]   io_out64_43,
  output [3:0]   io_out64_44,
  output [3:0]   io_out64_45,
  output [3:0]   io_out64_46,
  output [3:0]   io_out64_47,
  output [3:0]   io_out64_48,
  output [3:0]   io_out64_49,
  output [3:0]   io_out64_50,
  output [3:0]   io_out64_51,
  output [3:0]   io_out64_52,
  output [3:0]   io_out64_53,
  output [3:0]   io_out64_54,
  output [3:0]   io_out64_55,
  output [3:0]   io_out64_56,
  output [3:0]   io_out64_57,
  output [3:0]   io_out64_58,
  output [3:0]   io_out64_59,
  output [3:0]   io_out64_60,
  output [3:0]   io_out64_61,
  output [3:0]   io_out64_62,
  output [3:0]   io_out64_63,
  output         io_validout64_0,
  output         io_validout64_1,
  output         io_validout64_2,
  output         io_validout64_3,
  output         io_validout64_4,
  output         io_validout64_5,
  output         io_validout64_6,
  output         io_validout64_7,
  output         io_validout64_8,
  output         io_validout64_9,
  output         io_validout64_10,
  output         io_validout64_11,
  output         io_validout64_12,
  output         io_validout64_13,
  output         io_validout64_14,
  output         io_validout64_15,
  output         io_validout64_16,
  output         io_validout64_17,
  output         io_validout64_18,
  output         io_validout64_19,
  output         io_validout64_20,
  output         io_validout64_21,
  output         io_validout64_22,
  output         io_validout64_23,
  output         io_validout64_24,
  output         io_validout64_25,
  output         io_validout64_26,
  output         io_validout64_27,
  output         io_validout64_28,
  output         io_validout64_29,
  output         io_validout64_30,
  output         io_validout64_31,
  output         io_validout64_32,
  output         io_validout64_33,
  output         io_validout64_34,
  output         io_validout64_35,
  output         io_validout64_36,
  output         io_validout64_37,
  output         io_validout64_38,
  output         io_validout64_39,
  output         io_validout64_40,
  output         io_validout64_41,
  output         io_validout64_42,
  output         io_validout64_43,
  output         io_validout64_44,
  output         io_validout64_45,
  output         io_validout64_46,
  output         io_validout64_47,
  output         io_validout64_48,
  output         io_validout64_49,
  output         io_validout64_50,
  output         io_validout64_51,
  output         io_validout64_52,
  output         io_validout64_53,
  output         io_validout64_54,
  output         io_validout64_55,
  output         io_validout64_56,
  output         io_validout64_57,
  output         io_validout64_58,
  output         io_validout64_59,
  output         io_validout64_60,
  output         io_validout64_61,
  output         io_validout64_62,
  output         io_validout64_63,
  output [7:0]   io_addrout,
  input  [127:0] io_ctrl
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  egress2_0_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_0_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_0_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_1_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_1_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_1_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_2_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_2_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_2_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_3_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_3_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_3_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_4_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_4_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_4_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_5_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_5_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_5_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_6_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_6_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_6_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_7_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_7_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_7_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_8_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_8_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_8_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_9_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_9_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_9_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_10_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_10_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_10_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_11_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_11_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_11_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_12_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_12_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_12_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_13_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_13_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_13_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_14_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_14_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_14_io_ctrl; // @[BuildingBlock.scala 192:51]
  wire  egress2_15_clock; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_in4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_in4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_in4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_in4_3; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_out4_0; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_out4_1; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_out4_2; // @[BuildingBlock.scala 192:51]
  wire [4:0] egress2_15_io_out4_3; // @[BuildingBlock.scala 192:51]
  wire [7:0] egress2_15_io_ctrl; // @[BuildingBlock.scala 192:51]
  reg [7:0] addr; // @[BuildingBlock.scala 195:21]
  CLOScell4 egress2_0 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_0_clock),
    .io_in4_0(egress2_0_io_in4_0),
    .io_in4_1(egress2_0_io_in4_1),
    .io_in4_2(egress2_0_io_in4_2),
    .io_in4_3(egress2_0_io_in4_3),
    .io_out4_0(egress2_0_io_out4_0),
    .io_out4_1(egress2_0_io_out4_1),
    .io_out4_2(egress2_0_io_out4_2),
    .io_out4_3(egress2_0_io_out4_3),
    .io_ctrl(egress2_0_io_ctrl)
  );
  CLOScell4 egress2_1 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_1_clock),
    .io_in4_0(egress2_1_io_in4_0),
    .io_in4_1(egress2_1_io_in4_1),
    .io_in4_2(egress2_1_io_in4_2),
    .io_in4_3(egress2_1_io_in4_3),
    .io_out4_0(egress2_1_io_out4_0),
    .io_out4_1(egress2_1_io_out4_1),
    .io_out4_2(egress2_1_io_out4_2),
    .io_out4_3(egress2_1_io_out4_3),
    .io_ctrl(egress2_1_io_ctrl)
  );
  CLOScell4 egress2_2 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_2_clock),
    .io_in4_0(egress2_2_io_in4_0),
    .io_in4_1(egress2_2_io_in4_1),
    .io_in4_2(egress2_2_io_in4_2),
    .io_in4_3(egress2_2_io_in4_3),
    .io_out4_0(egress2_2_io_out4_0),
    .io_out4_1(egress2_2_io_out4_1),
    .io_out4_2(egress2_2_io_out4_2),
    .io_out4_3(egress2_2_io_out4_3),
    .io_ctrl(egress2_2_io_ctrl)
  );
  CLOScell4 egress2_3 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_3_clock),
    .io_in4_0(egress2_3_io_in4_0),
    .io_in4_1(egress2_3_io_in4_1),
    .io_in4_2(egress2_3_io_in4_2),
    .io_in4_3(egress2_3_io_in4_3),
    .io_out4_0(egress2_3_io_out4_0),
    .io_out4_1(egress2_3_io_out4_1),
    .io_out4_2(egress2_3_io_out4_2),
    .io_out4_3(egress2_3_io_out4_3),
    .io_ctrl(egress2_3_io_ctrl)
  );
  CLOScell4 egress2_4 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_4_clock),
    .io_in4_0(egress2_4_io_in4_0),
    .io_in4_1(egress2_4_io_in4_1),
    .io_in4_2(egress2_4_io_in4_2),
    .io_in4_3(egress2_4_io_in4_3),
    .io_out4_0(egress2_4_io_out4_0),
    .io_out4_1(egress2_4_io_out4_1),
    .io_out4_2(egress2_4_io_out4_2),
    .io_out4_3(egress2_4_io_out4_3),
    .io_ctrl(egress2_4_io_ctrl)
  );
  CLOScell4 egress2_5 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_5_clock),
    .io_in4_0(egress2_5_io_in4_0),
    .io_in4_1(egress2_5_io_in4_1),
    .io_in4_2(egress2_5_io_in4_2),
    .io_in4_3(egress2_5_io_in4_3),
    .io_out4_0(egress2_5_io_out4_0),
    .io_out4_1(egress2_5_io_out4_1),
    .io_out4_2(egress2_5_io_out4_2),
    .io_out4_3(egress2_5_io_out4_3),
    .io_ctrl(egress2_5_io_ctrl)
  );
  CLOScell4 egress2_6 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_6_clock),
    .io_in4_0(egress2_6_io_in4_0),
    .io_in4_1(egress2_6_io_in4_1),
    .io_in4_2(egress2_6_io_in4_2),
    .io_in4_3(egress2_6_io_in4_3),
    .io_out4_0(egress2_6_io_out4_0),
    .io_out4_1(egress2_6_io_out4_1),
    .io_out4_2(egress2_6_io_out4_2),
    .io_out4_3(egress2_6_io_out4_3),
    .io_ctrl(egress2_6_io_ctrl)
  );
  CLOScell4 egress2_7 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_7_clock),
    .io_in4_0(egress2_7_io_in4_0),
    .io_in4_1(egress2_7_io_in4_1),
    .io_in4_2(egress2_7_io_in4_2),
    .io_in4_3(egress2_7_io_in4_3),
    .io_out4_0(egress2_7_io_out4_0),
    .io_out4_1(egress2_7_io_out4_1),
    .io_out4_2(egress2_7_io_out4_2),
    .io_out4_3(egress2_7_io_out4_3),
    .io_ctrl(egress2_7_io_ctrl)
  );
  CLOScell4 egress2_8 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_8_clock),
    .io_in4_0(egress2_8_io_in4_0),
    .io_in4_1(egress2_8_io_in4_1),
    .io_in4_2(egress2_8_io_in4_2),
    .io_in4_3(egress2_8_io_in4_3),
    .io_out4_0(egress2_8_io_out4_0),
    .io_out4_1(egress2_8_io_out4_1),
    .io_out4_2(egress2_8_io_out4_2),
    .io_out4_3(egress2_8_io_out4_3),
    .io_ctrl(egress2_8_io_ctrl)
  );
  CLOScell4 egress2_9 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_9_clock),
    .io_in4_0(egress2_9_io_in4_0),
    .io_in4_1(egress2_9_io_in4_1),
    .io_in4_2(egress2_9_io_in4_2),
    .io_in4_3(egress2_9_io_in4_3),
    .io_out4_0(egress2_9_io_out4_0),
    .io_out4_1(egress2_9_io_out4_1),
    .io_out4_2(egress2_9_io_out4_2),
    .io_out4_3(egress2_9_io_out4_3),
    .io_ctrl(egress2_9_io_ctrl)
  );
  CLOScell4 egress2_10 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_10_clock),
    .io_in4_0(egress2_10_io_in4_0),
    .io_in4_1(egress2_10_io_in4_1),
    .io_in4_2(egress2_10_io_in4_2),
    .io_in4_3(egress2_10_io_in4_3),
    .io_out4_0(egress2_10_io_out4_0),
    .io_out4_1(egress2_10_io_out4_1),
    .io_out4_2(egress2_10_io_out4_2),
    .io_out4_3(egress2_10_io_out4_3),
    .io_ctrl(egress2_10_io_ctrl)
  );
  CLOScell4 egress2_11 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_11_clock),
    .io_in4_0(egress2_11_io_in4_0),
    .io_in4_1(egress2_11_io_in4_1),
    .io_in4_2(egress2_11_io_in4_2),
    .io_in4_3(egress2_11_io_in4_3),
    .io_out4_0(egress2_11_io_out4_0),
    .io_out4_1(egress2_11_io_out4_1),
    .io_out4_2(egress2_11_io_out4_2),
    .io_out4_3(egress2_11_io_out4_3),
    .io_ctrl(egress2_11_io_ctrl)
  );
  CLOScell4 egress2_12 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_12_clock),
    .io_in4_0(egress2_12_io_in4_0),
    .io_in4_1(egress2_12_io_in4_1),
    .io_in4_2(egress2_12_io_in4_2),
    .io_in4_3(egress2_12_io_in4_3),
    .io_out4_0(egress2_12_io_out4_0),
    .io_out4_1(egress2_12_io_out4_1),
    .io_out4_2(egress2_12_io_out4_2),
    .io_out4_3(egress2_12_io_out4_3),
    .io_ctrl(egress2_12_io_ctrl)
  );
  CLOScell4 egress2_13 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_13_clock),
    .io_in4_0(egress2_13_io_in4_0),
    .io_in4_1(egress2_13_io_in4_1),
    .io_in4_2(egress2_13_io_in4_2),
    .io_in4_3(egress2_13_io_in4_3),
    .io_out4_0(egress2_13_io_out4_0),
    .io_out4_1(egress2_13_io_out4_1),
    .io_out4_2(egress2_13_io_out4_2),
    .io_out4_3(egress2_13_io_out4_3),
    .io_ctrl(egress2_13_io_ctrl)
  );
  CLOScell4 egress2_14 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_14_clock),
    .io_in4_0(egress2_14_io_in4_0),
    .io_in4_1(egress2_14_io_in4_1),
    .io_in4_2(egress2_14_io_in4_2),
    .io_in4_3(egress2_14_io_in4_3),
    .io_out4_0(egress2_14_io_out4_0),
    .io_out4_1(egress2_14_io_out4_1),
    .io_out4_2(egress2_14_io_out4_2),
    .io_out4_3(egress2_14_io_out4_3),
    .io_ctrl(egress2_14_io_ctrl)
  );
  CLOScell4 egress2_15 ( // @[BuildingBlock.scala 192:51]
    .clock(egress2_15_clock),
    .io_in4_0(egress2_15_io_in4_0),
    .io_in4_1(egress2_15_io_in4_1),
    .io_in4_2(egress2_15_io_in4_2),
    .io_in4_3(egress2_15_io_in4_3),
    .io_out4_0(egress2_15_io_out4_0),
    .io_out4_1(egress2_15_io_out4_1),
    .io_out4_2(egress2_15_io_out4_2),
    .io_out4_3(egress2_15_io_out4_3),
    .io_ctrl(egress2_15_io_ctrl)
  );
  assign io_out64_0 = egress2_0_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_1 = egress2_0_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_2 = egress2_0_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_3 = egress2_0_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_4 = egress2_1_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_5 = egress2_1_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_6 = egress2_1_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_7 = egress2_1_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_8 = egress2_2_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_9 = egress2_2_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_10 = egress2_2_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_11 = egress2_2_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_12 = egress2_3_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_13 = egress2_3_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_14 = egress2_3_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_15 = egress2_3_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_16 = egress2_4_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_17 = egress2_4_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_18 = egress2_4_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_19 = egress2_4_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_20 = egress2_5_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_21 = egress2_5_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_22 = egress2_5_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_23 = egress2_5_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_24 = egress2_6_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_25 = egress2_6_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_26 = egress2_6_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_27 = egress2_6_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_28 = egress2_7_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_29 = egress2_7_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_30 = egress2_7_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_31 = egress2_7_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_32 = egress2_8_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_33 = egress2_8_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_34 = egress2_8_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_35 = egress2_8_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_36 = egress2_9_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_37 = egress2_9_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_38 = egress2_9_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_39 = egress2_9_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_40 = egress2_10_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_41 = egress2_10_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_42 = egress2_10_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_43 = egress2_10_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_44 = egress2_11_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_45 = egress2_11_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_46 = egress2_11_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_47 = egress2_11_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_48 = egress2_12_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_49 = egress2_12_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_50 = egress2_12_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_51 = egress2_12_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_52 = egress2_13_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_53 = egress2_13_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_54 = egress2_13_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_55 = egress2_13_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_56 = egress2_14_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_57 = egress2_14_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_58 = egress2_14_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_59 = egress2_14_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_60 = egress2_15_io_out4_0[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_61 = egress2_15_io_out4_1[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_62 = egress2_15_io_out4_2[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_out64_63 = egress2_15_io_out4_3[3:0]; // @[BuildingBlock.scala 206:47]
  assign io_validout64_0 = egress2_0_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_1 = egress2_0_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_2 = egress2_0_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_3 = egress2_0_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_4 = egress2_1_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_5 = egress2_1_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_6 = egress2_1_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_7 = egress2_1_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_8 = egress2_2_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_9 = egress2_2_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_10 = egress2_2_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_11 = egress2_2_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_12 = egress2_3_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_13 = egress2_3_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_14 = egress2_3_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_15 = egress2_3_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_16 = egress2_4_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_17 = egress2_4_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_18 = egress2_4_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_19 = egress2_4_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_20 = egress2_5_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_21 = egress2_5_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_22 = egress2_5_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_23 = egress2_5_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_24 = egress2_6_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_25 = egress2_6_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_26 = egress2_6_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_27 = egress2_6_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_28 = egress2_7_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_29 = egress2_7_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_30 = egress2_7_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_31 = egress2_7_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_32 = egress2_8_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_33 = egress2_8_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_34 = egress2_8_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_35 = egress2_8_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_36 = egress2_9_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_37 = egress2_9_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_38 = egress2_9_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_39 = egress2_9_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_40 = egress2_10_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_41 = egress2_10_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_42 = egress2_10_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_43 = egress2_10_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_44 = egress2_11_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_45 = egress2_11_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_46 = egress2_11_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_47 = egress2_11_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_48 = egress2_12_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_49 = egress2_12_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_50 = egress2_12_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_51 = egress2_12_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_52 = egress2_13_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_53 = egress2_13_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_54 = egress2_13_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_55 = egress2_13_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_56 = egress2_14_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_57 = egress2_14_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_58 = egress2_14_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_59 = egress2_14_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_60 = egress2_15_io_out4_0[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_61 = egress2_15_io_out4_1[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_62 = egress2_15_io_out4_2[4]; // @[BuildingBlock.scala 207:52]
  assign io_validout64_63 = egress2_15_io_out4_3[4]; // @[BuildingBlock.scala 207:52]
  assign io_addrout = addr; // @[BuildingBlock.scala 196:14]
  assign egress2_0_clock = clock;
  assign egress2_0_io_in4_0 = {io_validin64_0,io_in64_0}; // @[Cat.scala 30:58]
  assign egress2_0_io_in4_1 = {io_validin64_1,io_in64_1}; // @[Cat.scala 30:58]
  assign egress2_0_io_in4_2 = {io_validin64_2,io_in64_2}; // @[Cat.scala 30:58]
  assign egress2_0_io_in4_3 = {io_validin64_3,io_in64_3}; // @[Cat.scala 30:58]
  assign egress2_0_io_ctrl = io_ctrl[127:120]; // @[BuildingBlock.scala 211:34]
  assign egress2_1_clock = clock;
  assign egress2_1_io_in4_0 = {io_validin64_4,io_in64_4}; // @[Cat.scala 30:58]
  assign egress2_1_io_in4_1 = {io_validin64_5,io_in64_5}; // @[Cat.scala 30:58]
  assign egress2_1_io_in4_2 = {io_validin64_6,io_in64_6}; // @[Cat.scala 30:58]
  assign egress2_1_io_in4_3 = {io_validin64_7,io_in64_7}; // @[Cat.scala 30:58]
  assign egress2_1_io_ctrl = io_ctrl[119:112]; // @[BuildingBlock.scala 211:34]
  assign egress2_2_clock = clock;
  assign egress2_2_io_in4_0 = {io_validin64_8,io_in64_8}; // @[Cat.scala 30:58]
  assign egress2_2_io_in4_1 = {io_validin64_9,io_in64_9}; // @[Cat.scala 30:58]
  assign egress2_2_io_in4_2 = {io_validin64_10,io_in64_10}; // @[Cat.scala 30:58]
  assign egress2_2_io_in4_3 = {io_validin64_11,io_in64_11}; // @[Cat.scala 30:58]
  assign egress2_2_io_ctrl = io_ctrl[111:104]; // @[BuildingBlock.scala 211:34]
  assign egress2_3_clock = clock;
  assign egress2_3_io_in4_0 = {io_validin64_12,io_in64_12}; // @[Cat.scala 30:58]
  assign egress2_3_io_in4_1 = {io_validin64_13,io_in64_13}; // @[Cat.scala 30:58]
  assign egress2_3_io_in4_2 = {io_validin64_14,io_in64_14}; // @[Cat.scala 30:58]
  assign egress2_3_io_in4_3 = {io_validin64_15,io_in64_15}; // @[Cat.scala 30:58]
  assign egress2_3_io_ctrl = io_ctrl[103:96]; // @[BuildingBlock.scala 211:34]
  assign egress2_4_clock = clock;
  assign egress2_4_io_in4_0 = {io_validin64_16,io_in64_16}; // @[Cat.scala 30:58]
  assign egress2_4_io_in4_1 = {io_validin64_17,io_in64_17}; // @[Cat.scala 30:58]
  assign egress2_4_io_in4_2 = {io_validin64_18,io_in64_18}; // @[Cat.scala 30:58]
  assign egress2_4_io_in4_3 = {io_validin64_19,io_in64_19}; // @[Cat.scala 30:58]
  assign egress2_4_io_ctrl = io_ctrl[95:88]; // @[BuildingBlock.scala 211:34]
  assign egress2_5_clock = clock;
  assign egress2_5_io_in4_0 = {io_validin64_20,io_in64_20}; // @[Cat.scala 30:58]
  assign egress2_5_io_in4_1 = {io_validin64_21,io_in64_21}; // @[Cat.scala 30:58]
  assign egress2_5_io_in4_2 = {io_validin64_22,io_in64_22}; // @[Cat.scala 30:58]
  assign egress2_5_io_in4_3 = {io_validin64_23,io_in64_23}; // @[Cat.scala 30:58]
  assign egress2_5_io_ctrl = io_ctrl[87:80]; // @[BuildingBlock.scala 211:34]
  assign egress2_6_clock = clock;
  assign egress2_6_io_in4_0 = {io_validin64_24,io_in64_24}; // @[Cat.scala 30:58]
  assign egress2_6_io_in4_1 = {io_validin64_25,io_in64_25}; // @[Cat.scala 30:58]
  assign egress2_6_io_in4_2 = {io_validin64_26,io_in64_26}; // @[Cat.scala 30:58]
  assign egress2_6_io_in4_3 = {io_validin64_27,io_in64_27}; // @[Cat.scala 30:58]
  assign egress2_6_io_ctrl = io_ctrl[79:72]; // @[BuildingBlock.scala 211:34]
  assign egress2_7_clock = clock;
  assign egress2_7_io_in4_0 = {io_validin64_28,io_in64_28}; // @[Cat.scala 30:58]
  assign egress2_7_io_in4_1 = {io_validin64_29,io_in64_29}; // @[Cat.scala 30:58]
  assign egress2_7_io_in4_2 = {io_validin64_30,io_in64_30}; // @[Cat.scala 30:58]
  assign egress2_7_io_in4_3 = {io_validin64_31,io_in64_31}; // @[Cat.scala 30:58]
  assign egress2_7_io_ctrl = io_ctrl[71:64]; // @[BuildingBlock.scala 211:34]
  assign egress2_8_clock = clock;
  assign egress2_8_io_in4_0 = {io_validin64_32,io_in64_32}; // @[Cat.scala 30:58]
  assign egress2_8_io_in4_1 = {io_validin64_33,io_in64_33}; // @[Cat.scala 30:58]
  assign egress2_8_io_in4_2 = {io_validin64_34,io_in64_34}; // @[Cat.scala 30:58]
  assign egress2_8_io_in4_3 = {io_validin64_35,io_in64_35}; // @[Cat.scala 30:58]
  assign egress2_8_io_ctrl = io_ctrl[63:56]; // @[BuildingBlock.scala 211:34]
  assign egress2_9_clock = clock;
  assign egress2_9_io_in4_0 = {io_validin64_36,io_in64_36}; // @[Cat.scala 30:58]
  assign egress2_9_io_in4_1 = {io_validin64_37,io_in64_37}; // @[Cat.scala 30:58]
  assign egress2_9_io_in4_2 = {io_validin64_38,io_in64_38}; // @[Cat.scala 30:58]
  assign egress2_9_io_in4_3 = {io_validin64_39,io_in64_39}; // @[Cat.scala 30:58]
  assign egress2_9_io_ctrl = io_ctrl[55:48]; // @[BuildingBlock.scala 211:34]
  assign egress2_10_clock = clock;
  assign egress2_10_io_in4_0 = {io_validin64_40,io_in64_40}; // @[Cat.scala 30:58]
  assign egress2_10_io_in4_1 = {io_validin64_41,io_in64_41}; // @[Cat.scala 30:58]
  assign egress2_10_io_in4_2 = {io_validin64_42,io_in64_42}; // @[Cat.scala 30:58]
  assign egress2_10_io_in4_3 = {io_validin64_43,io_in64_43}; // @[Cat.scala 30:58]
  assign egress2_10_io_ctrl = io_ctrl[47:40]; // @[BuildingBlock.scala 211:34]
  assign egress2_11_clock = clock;
  assign egress2_11_io_in4_0 = {io_validin64_44,io_in64_44}; // @[Cat.scala 30:58]
  assign egress2_11_io_in4_1 = {io_validin64_45,io_in64_45}; // @[Cat.scala 30:58]
  assign egress2_11_io_in4_2 = {io_validin64_46,io_in64_46}; // @[Cat.scala 30:58]
  assign egress2_11_io_in4_3 = {io_validin64_47,io_in64_47}; // @[Cat.scala 30:58]
  assign egress2_11_io_ctrl = io_ctrl[39:32]; // @[BuildingBlock.scala 211:34]
  assign egress2_12_clock = clock;
  assign egress2_12_io_in4_0 = {io_validin64_48,io_in64_48}; // @[Cat.scala 30:58]
  assign egress2_12_io_in4_1 = {io_validin64_49,io_in64_49}; // @[Cat.scala 30:58]
  assign egress2_12_io_in4_2 = {io_validin64_50,io_in64_50}; // @[Cat.scala 30:58]
  assign egress2_12_io_in4_3 = {io_validin64_51,io_in64_51}; // @[Cat.scala 30:58]
  assign egress2_12_io_ctrl = io_ctrl[31:24]; // @[BuildingBlock.scala 211:34]
  assign egress2_13_clock = clock;
  assign egress2_13_io_in4_0 = {io_validin64_52,io_in64_52}; // @[Cat.scala 30:58]
  assign egress2_13_io_in4_1 = {io_validin64_53,io_in64_53}; // @[Cat.scala 30:58]
  assign egress2_13_io_in4_2 = {io_validin64_54,io_in64_54}; // @[Cat.scala 30:58]
  assign egress2_13_io_in4_3 = {io_validin64_55,io_in64_55}; // @[Cat.scala 30:58]
  assign egress2_13_io_ctrl = io_ctrl[23:16]; // @[BuildingBlock.scala 211:34]
  assign egress2_14_clock = clock;
  assign egress2_14_io_in4_0 = {io_validin64_56,io_in64_56}; // @[Cat.scala 30:58]
  assign egress2_14_io_in4_1 = {io_validin64_57,io_in64_57}; // @[Cat.scala 30:58]
  assign egress2_14_io_in4_2 = {io_validin64_58,io_in64_58}; // @[Cat.scala 30:58]
  assign egress2_14_io_in4_3 = {io_validin64_59,io_in64_59}; // @[Cat.scala 30:58]
  assign egress2_14_io_ctrl = io_ctrl[15:8]; // @[BuildingBlock.scala 211:34]
  assign egress2_15_clock = clock;
  assign egress2_15_io_in4_0 = {io_validin64_60,io_in64_60}; // @[Cat.scala 30:58]
  assign egress2_15_io_in4_1 = {io_validin64_61,io_in64_61}; // @[Cat.scala 30:58]
  assign egress2_15_io_in4_2 = {io_validin64_62,io_in64_62}; // @[Cat.scala 30:58]
  assign egress2_15_io_in4_3 = {io_validin64_63,io_in64_63}; // @[Cat.scala 30:58]
  assign egress2_15_io_ctrl = io_ctrl[7:0]; // @[BuildingBlock.scala 211:34]
  always @(posedge clock) begin
    addr <= io_addrin; // @[BuildingBlock.scala 195:21]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  addr = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BuildingBlockNew(
  input          clock,
  input          reset,
  input  [3:0]   io_d_in_0_a,
  input          io_d_in_0_valid_a,
  input  [3:0]   io_d_in_0_b,
  input          io_d_in_0_valid_b,
  input  [3:0]   io_d_in_1_a,
  input          io_d_in_1_valid_a,
  input  [3:0]   io_d_in_1_b,
  input          io_d_in_1_valid_b,
  input  [3:0]   io_d_in_2_a,
  input          io_d_in_2_valid_a,
  input  [3:0]   io_d_in_2_b,
  input          io_d_in_2_valid_b,
  input  [3:0]   io_d_in_3_a,
  input          io_d_in_3_valid_a,
  input  [3:0]   io_d_in_3_b,
  input          io_d_in_3_valid_b,
  input  [3:0]   io_d_in_4_a,
  input          io_d_in_4_valid_a,
  input  [3:0]   io_d_in_4_b,
  input          io_d_in_4_valid_b,
  input  [3:0]   io_d_in_5_a,
  input          io_d_in_5_valid_a,
  input  [3:0]   io_d_in_5_b,
  input          io_d_in_5_valid_b,
  input  [3:0]   io_d_in_6_a,
  input          io_d_in_6_valid_a,
  input  [3:0]   io_d_in_6_b,
  input          io_d_in_6_valid_b,
  input  [3:0]   io_d_in_7_a,
  input          io_d_in_7_valid_a,
  input  [3:0]   io_d_in_7_b,
  input          io_d_in_7_valid_b,
  input  [3:0]   io_d_in_8_a,
  input          io_d_in_8_valid_a,
  input  [3:0]   io_d_in_8_b,
  input          io_d_in_8_valid_b,
  input  [3:0]   io_d_in_9_a,
  input          io_d_in_9_valid_a,
  input  [3:0]   io_d_in_9_b,
  input          io_d_in_9_valid_b,
  input  [3:0]   io_d_in_10_a,
  input          io_d_in_10_valid_a,
  input  [3:0]   io_d_in_10_b,
  input          io_d_in_10_valid_b,
  input  [3:0]   io_d_in_11_a,
  input          io_d_in_11_valid_a,
  input  [3:0]   io_d_in_11_b,
  input          io_d_in_11_valid_b,
  input  [3:0]   io_d_in_12_a,
  input          io_d_in_12_valid_a,
  input  [3:0]   io_d_in_12_b,
  input          io_d_in_12_valid_b,
  input  [3:0]   io_d_in_13_a,
  input          io_d_in_13_valid_a,
  input  [3:0]   io_d_in_13_b,
  input          io_d_in_13_valid_b,
  input  [3:0]   io_d_in_14_a,
  input          io_d_in_14_valid_a,
  input  [3:0]   io_d_in_14_b,
  input          io_d_in_14_valid_b,
  input  [3:0]   io_d_in_15_a,
  input          io_d_in_15_valid_a,
  input  [3:0]   io_d_in_15_b,
  input          io_d_in_15_valid_b,
  input  [3:0]   io_d_in_16_a,
  input          io_d_in_16_valid_a,
  input  [3:0]   io_d_in_16_b,
  input          io_d_in_16_valid_b,
  input  [3:0]   io_d_in_17_a,
  input          io_d_in_17_valid_a,
  input  [3:0]   io_d_in_17_b,
  input          io_d_in_17_valid_b,
  input  [3:0]   io_d_in_18_a,
  input          io_d_in_18_valid_a,
  input  [3:0]   io_d_in_18_b,
  input          io_d_in_18_valid_b,
  input  [3:0]   io_d_in_19_a,
  input          io_d_in_19_valid_a,
  input  [3:0]   io_d_in_19_b,
  input          io_d_in_19_valid_b,
  input  [3:0]   io_d_in_20_a,
  input          io_d_in_20_valid_a,
  input  [3:0]   io_d_in_20_b,
  input          io_d_in_20_valid_b,
  input  [3:0]   io_d_in_21_a,
  input          io_d_in_21_valid_a,
  input  [3:0]   io_d_in_21_b,
  input          io_d_in_21_valid_b,
  input  [3:0]   io_d_in_22_a,
  input          io_d_in_22_valid_a,
  input  [3:0]   io_d_in_22_b,
  input          io_d_in_22_valid_b,
  input  [3:0]   io_d_in_23_a,
  input          io_d_in_23_valid_a,
  input  [3:0]   io_d_in_23_b,
  input          io_d_in_23_valid_b,
  input  [3:0]   io_d_in_24_a,
  input          io_d_in_24_valid_a,
  input  [3:0]   io_d_in_24_b,
  input          io_d_in_24_valid_b,
  input  [3:0]   io_d_in_25_a,
  input          io_d_in_25_valid_a,
  input  [3:0]   io_d_in_25_b,
  input          io_d_in_25_valid_b,
  input  [3:0]   io_d_in_26_a,
  input          io_d_in_26_valid_a,
  input  [3:0]   io_d_in_26_b,
  input          io_d_in_26_valid_b,
  input  [3:0]   io_d_in_27_a,
  input          io_d_in_27_valid_a,
  input  [3:0]   io_d_in_27_b,
  input          io_d_in_27_valid_b,
  input  [3:0]   io_d_in_28_a,
  input          io_d_in_28_valid_a,
  input  [3:0]   io_d_in_28_b,
  input          io_d_in_28_valid_b,
  input  [3:0]   io_d_in_29_a,
  input          io_d_in_29_valid_a,
  input  [3:0]   io_d_in_29_b,
  input          io_d_in_29_valid_b,
  input  [3:0]   io_d_in_30_a,
  input          io_d_in_30_valid_a,
  input  [3:0]   io_d_in_30_b,
  input          io_d_in_30_valid_b,
  input  [3:0]   io_d_in_31_a,
  input          io_d_in_31_valid_a,
  input  [3:0]   io_d_in_31_b,
  input          io_d_in_31_valid_b,
  output [3:0]   io_d_out_0_a,
  output         io_d_out_0_valid_a,
  output [3:0]   io_d_out_0_b,
  output         io_d_out_0_valid_b,
  output [3:0]   io_d_out_1_a,
  output         io_d_out_1_valid_a,
  output [3:0]   io_d_out_1_b,
  output         io_d_out_1_valid_b,
  output [3:0]   io_d_out_2_a,
  output         io_d_out_2_valid_a,
  output [3:0]   io_d_out_2_b,
  output         io_d_out_2_valid_b,
  output [3:0]   io_d_out_3_a,
  output         io_d_out_3_valid_a,
  output [3:0]   io_d_out_3_b,
  output         io_d_out_3_valid_b,
  output [3:0]   io_d_out_4_a,
  output         io_d_out_4_valid_a,
  output [3:0]   io_d_out_4_b,
  output         io_d_out_4_valid_b,
  output [3:0]   io_d_out_5_a,
  output         io_d_out_5_valid_a,
  output [3:0]   io_d_out_5_b,
  output         io_d_out_5_valid_b,
  output [3:0]   io_d_out_6_a,
  output         io_d_out_6_valid_a,
  output [3:0]   io_d_out_6_b,
  output         io_d_out_6_valid_b,
  output [3:0]   io_d_out_7_a,
  output         io_d_out_7_valid_a,
  output [3:0]   io_d_out_7_b,
  output         io_d_out_7_valid_b,
  output [3:0]   io_d_out_8_a,
  output         io_d_out_8_valid_a,
  output [3:0]   io_d_out_8_b,
  output         io_d_out_8_valid_b,
  output [3:0]   io_d_out_9_a,
  output         io_d_out_9_valid_a,
  output [3:0]   io_d_out_9_b,
  output         io_d_out_9_valid_b,
  output [3:0]   io_d_out_10_a,
  output         io_d_out_10_valid_a,
  output [3:0]   io_d_out_10_b,
  output         io_d_out_10_valid_b,
  output [3:0]   io_d_out_11_a,
  output         io_d_out_11_valid_a,
  output [3:0]   io_d_out_11_b,
  output         io_d_out_11_valid_b,
  output [3:0]   io_d_out_12_a,
  output         io_d_out_12_valid_a,
  output [3:0]   io_d_out_12_b,
  output         io_d_out_12_valid_b,
  output [3:0]   io_d_out_13_a,
  output         io_d_out_13_valid_a,
  output [3:0]   io_d_out_13_b,
  output         io_d_out_13_valid_b,
  output [3:0]   io_d_out_14_a,
  output         io_d_out_14_valid_a,
  output [3:0]   io_d_out_14_b,
  output         io_d_out_14_valid_b,
  output [3:0]   io_d_out_15_a,
  output         io_d_out_15_valid_a,
  output [3:0]   io_d_out_15_b,
  output         io_d_out_15_valid_b,
  output [3:0]   io_d_out_16_a,
  output         io_d_out_16_valid_a,
  output [3:0]   io_d_out_16_b,
  output         io_d_out_16_valid_b,
  output [3:0]   io_d_out_17_a,
  output         io_d_out_17_valid_a,
  output [3:0]   io_d_out_17_b,
  output         io_d_out_17_valid_b,
  output [3:0]   io_d_out_18_a,
  output         io_d_out_18_valid_a,
  output [3:0]   io_d_out_18_b,
  output         io_d_out_18_valid_b,
  output [3:0]   io_d_out_19_a,
  output         io_d_out_19_valid_a,
  output [3:0]   io_d_out_19_b,
  output         io_d_out_19_valid_b,
  output [3:0]   io_d_out_20_a,
  output         io_d_out_20_valid_a,
  output [3:0]   io_d_out_20_b,
  output         io_d_out_20_valid_b,
  output [3:0]   io_d_out_21_a,
  output         io_d_out_21_valid_a,
  output [3:0]   io_d_out_21_b,
  output         io_d_out_21_valid_b,
  output [3:0]   io_d_out_22_a,
  output         io_d_out_22_valid_a,
  output [3:0]   io_d_out_22_b,
  output         io_d_out_22_valid_b,
  output [3:0]   io_d_out_23_a,
  output         io_d_out_23_valid_a,
  output [3:0]   io_d_out_23_b,
  output         io_d_out_23_valid_b,
  output [3:0]   io_d_out_24_a,
  output         io_d_out_24_valid_a,
  output [3:0]   io_d_out_24_b,
  output         io_d_out_24_valid_b,
  output [3:0]   io_d_out_25_a,
  output         io_d_out_25_valid_a,
  output [3:0]   io_d_out_25_b,
  output         io_d_out_25_valid_b,
  output [3:0]   io_d_out_26_a,
  output         io_d_out_26_valid_a,
  output [3:0]   io_d_out_26_b,
  output         io_d_out_26_valid_b,
  output [3:0]   io_d_out_27_a,
  output         io_d_out_27_valid_a,
  output [3:0]   io_d_out_27_b,
  output         io_d_out_27_valid_b,
  output [3:0]   io_d_out_28_a,
  output         io_d_out_28_valid_a,
  output [3:0]   io_d_out_28_b,
  output         io_d_out_28_valid_b,
  output [3:0]   io_d_out_29_a,
  output         io_d_out_29_valid_a,
  output [3:0]   io_d_out_29_b,
  output         io_d_out_29_valid_b,
  output [3:0]   io_d_out_30_a,
  output         io_d_out_30_valid_a,
  output [3:0]   io_d_out_30_b,
  output         io_d_out_30_valid_b,
  output [3:0]   io_d_out_31_a,
  output         io_d_out_31_valid_a,
  output [3:0]   io_d_out_31_b,
  output         io_d_out_31_valid_b,
  input          io_wr_en_mem1,
  input          io_wr_en_mem2,
  input          io_wr_en_mem3,
  input          io_wr_en_mem4,
  input          io_wr_en_mem5,
  input          io_wr_en_mem6,
  input  [287:0] io_wr_instr_mem1,
  input  [127:0] io_wr_instr_mem2,
  input  [127:0] io_wr_instr_mem3,
  input  [127:0] io_wr_instr_mem4,
  input  [127:0] io_wr_instr_mem5,
  input  [127:0] io_wr_instr_mem6,
  input  [7:0]   io_PC1_in,
  output [7:0]   io_PC6_out,
  input  [7:0]   io_Addr_in,
  output [7:0]   io_Addr_out
);
`ifdef RANDOMIZE_MEM_INIT
  reg [287:0] _RAND_0;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_4;
  reg [127:0] _RAND_6;
  reg [127:0] _RAND_8;
  reg [127:0] _RAND_10;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
`endif // RANDOMIZE_REG_INIT
  reg [287:0] Mem1 [0:255]; // @[BuildingBlockNew.scala 33:25]
  wire [287:0] Mem1_instr1_MPORT_data; // @[BuildingBlockNew.scala 33:25]
  wire [7:0] Mem1_instr1_MPORT_addr; // @[BuildingBlockNew.scala 33:25]
  wire [287:0] Mem1_MPORT_data; // @[BuildingBlockNew.scala 33:25]
  wire [7:0] Mem1_MPORT_addr; // @[BuildingBlockNew.scala 33:25]
  wire  Mem1_MPORT_mask; // @[BuildingBlockNew.scala 33:25]
  wire  Mem1_MPORT_en; // @[BuildingBlockNew.scala 33:25]
  reg [7:0] Mem1_instr1_MPORT_addr_pipe_0;
  reg [127:0] Mem2 [0:255]; // @[BuildingBlockNew.scala 34:25]
  wire [127:0] Mem2_instr2_MPORT_data; // @[BuildingBlockNew.scala 34:25]
  wire [7:0] Mem2_instr2_MPORT_addr; // @[BuildingBlockNew.scala 34:25]
  wire [127:0] Mem2_MPORT_1_data; // @[BuildingBlockNew.scala 34:25]
  wire [7:0] Mem2_MPORT_1_addr; // @[BuildingBlockNew.scala 34:25]
  wire  Mem2_MPORT_1_mask; // @[BuildingBlockNew.scala 34:25]
  wire  Mem2_MPORT_1_en; // @[BuildingBlockNew.scala 34:25]
  reg [7:0] Mem2_instr2_MPORT_addr_pipe_0;
  reg [127:0] Mem3 [0:255]; // @[BuildingBlockNew.scala 35:25]
  wire [127:0] Mem3_instr3_MPORT_data; // @[BuildingBlockNew.scala 35:25]
  wire [7:0] Mem3_instr3_MPORT_addr; // @[BuildingBlockNew.scala 35:25]
  wire [127:0] Mem3_MPORT_2_data; // @[BuildingBlockNew.scala 35:25]
  wire [7:0] Mem3_MPORT_2_addr; // @[BuildingBlockNew.scala 35:25]
  wire  Mem3_MPORT_2_mask; // @[BuildingBlockNew.scala 35:25]
  wire  Mem3_MPORT_2_en; // @[BuildingBlockNew.scala 35:25]
  reg [7:0] Mem3_instr3_MPORT_addr_pipe_0;
  reg [127:0] Mem4 [0:255]; // @[BuildingBlockNew.scala 36:25]
  wire [127:0] Mem4_instr4_MPORT_data; // @[BuildingBlockNew.scala 36:25]
  wire [7:0] Mem4_instr4_MPORT_addr; // @[BuildingBlockNew.scala 36:25]
  wire [127:0] Mem4_MPORT_3_data; // @[BuildingBlockNew.scala 36:25]
  wire [7:0] Mem4_MPORT_3_addr; // @[BuildingBlockNew.scala 36:25]
  wire  Mem4_MPORT_3_mask; // @[BuildingBlockNew.scala 36:25]
  wire  Mem4_MPORT_3_en; // @[BuildingBlockNew.scala 36:25]
  reg [7:0] Mem4_instr4_MPORT_addr_pipe_0;
  reg [127:0] Mem5 [0:255]; // @[BuildingBlockNew.scala 37:25]
  wire [127:0] Mem5_instr5_MPORT_data; // @[BuildingBlockNew.scala 37:25]
  wire [7:0] Mem5_instr5_MPORT_addr; // @[BuildingBlockNew.scala 37:25]
  wire [127:0] Mem5_MPORT_4_data; // @[BuildingBlockNew.scala 37:25]
  wire [7:0] Mem5_MPORT_4_addr; // @[BuildingBlockNew.scala 37:25]
  wire  Mem5_MPORT_4_mask; // @[BuildingBlockNew.scala 37:25]
  wire  Mem5_MPORT_4_en; // @[BuildingBlockNew.scala 37:25]
  reg [7:0] Mem5_instr5_MPORT_addr_pipe_0;
  reg [127:0] Mem6 [0:255]; // @[BuildingBlockNew.scala 38:25]
  wire [127:0] Mem6_instr6_MPORT_data; // @[BuildingBlockNew.scala 38:25]
  wire [7:0] Mem6_instr6_MPORT_addr; // @[BuildingBlockNew.scala 38:25]
  wire [127:0] Mem6_MPORT_5_data; // @[BuildingBlockNew.scala 38:25]
  wire [7:0] Mem6_MPORT_5_addr; // @[BuildingBlockNew.scala 38:25]
  wire  Mem6_MPORT_5_mask; // @[BuildingBlockNew.scala 38:25]
  wire  Mem6_MPORT_5_en; // @[BuildingBlockNew.scala 38:25]
  reg [7:0] Mem6_instr6_MPORT_addr_pipe_0;
  wire  peCol_clock; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_reset; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_0_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_0_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_0_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_0_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_1_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_1_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_1_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_1_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_2_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_2_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_2_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_2_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_3_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_3_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_3_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_3_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_4_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_4_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_4_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_4_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_5_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_5_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_5_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_5_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_6_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_6_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_6_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_6_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_7_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_7_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_7_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_7_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_8_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_8_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_8_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_8_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_9_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_9_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_9_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_9_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_10_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_10_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_10_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_10_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_11_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_11_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_11_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_11_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_12_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_12_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_12_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_12_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_13_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_13_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_13_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_13_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_14_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_14_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_14_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_14_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_15_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_15_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_15_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_15_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_16_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_16_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_16_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_16_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_17_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_17_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_17_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_17_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_18_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_18_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_18_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_18_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_19_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_19_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_19_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_19_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_20_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_20_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_20_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_20_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_21_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_21_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_21_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_21_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_22_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_22_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_22_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_22_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_23_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_23_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_23_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_23_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_24_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_24_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_24_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_24_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_25_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_25_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_25_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_25_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_26_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_26_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_26_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_26_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_27_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_27_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_27_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_27_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_28_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_28_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_28_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_28_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_29_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_29_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_29_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_29_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_30_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_30_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_30_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_30_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_31_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_31_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_in_31_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_in_31_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_0_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_0_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_0_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_0_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_1_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_1_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_1_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_1_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_2_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_2_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_2_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_2_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_3_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_3_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_3_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_3_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_4_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_4_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_4_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_4_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_5_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_5_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_5_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_5_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_6_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_6_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_6_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_6_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_7_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_7_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_7_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_7_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_8_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_8_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_8_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_8_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_9_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_9_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_9_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_9_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_10_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_10_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_10_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_10_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_11_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_11_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_11_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_11_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_12_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_12_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_12_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_12_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_13_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_13_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_13_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_13_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_14_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_14_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_14_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_14_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_15_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_15_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_15_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_15_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_16_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_16_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_16_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_16_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_17_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_17_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_17_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_17_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_18_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_18_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_18_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_18_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_19_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_19_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_19_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_19_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_20_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_20_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_20_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_20_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_21_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_21_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_21_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_21_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_22_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_22_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_22_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_22_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_23_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_23_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_23_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_23_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_24_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_24_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_24_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_24_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_25_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_25_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_25_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_25_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_26_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_26_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_26_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_26_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_27_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_27_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_27_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_27_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_28_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_28_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_28_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_28_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_29_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_29_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_29_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_29_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_30_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_30_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_30_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_30_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_31_a; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_31_valid_a; // @[BuildingBlockNew.scala 83:21]
  wire [3:0] peCol_io_d_out_31_b; // @[BuildingBlockNew.scala 83:21]
  wire  peCol_io_d_out_31_valid_b; // @[BuildingBlockNew.scala 83:21]
  wire [7:0] peCol_io_addrin; // @[BuildingBlockNew.scala 83:21]
  wire [7:0] peCol_io_addrout; // @[BuildingBlockNew.scala 83:21]
  wire [287:0] peCol_io_instr; // @[BuildingBlockNew.scala 83:21]
  wire  ingress1_clock; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_0; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_1; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_2; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_3; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_4; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_5; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_6; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_7; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_8; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_9; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_10; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_11; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_12; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_13; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_14; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_15; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_16; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_17; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_18; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_19; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_20; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_21; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_22; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_23; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_24; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_25; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_26; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_27; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_28; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_29; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_30; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_31; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_32; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_33; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_34; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_35; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_36; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_37; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_38; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_39; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_40; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_41; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_42; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_43; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_44; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_45; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_46; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_47; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_48; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_49; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_50; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_51; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_52; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_53; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_54; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_55; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_56; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_57; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_58; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_59; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_60; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_61; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_62; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_in64_63; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_0; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_1; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_2; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_3; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_4; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_5; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_6; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_7; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_8; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_9; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_10; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_11; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_12; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_13; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_14; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_15; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_16; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_17; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_18; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_19; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_20; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_21; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_22; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_23; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_24; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_25; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_26; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_27; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_28; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_29; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_30; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_31; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_32; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_33; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_34; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_35; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_36; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_37; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_38; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_39; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_40; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_41; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_42; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_43; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_44; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_45; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_46; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_47; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_48; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_49; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_50; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_51; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_52; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_53; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_54; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_55; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_56; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_57; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_58; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_59; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_60; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_61; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_62; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validin64_63; // @[BuildingBlockNew.scala 84:24]
  wire [7:0] ingress1_io_addrin; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_0; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_1; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_2; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_3; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_4; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_5; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_6; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_7; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_8; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_9; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_10; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_11; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_12; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_13; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_14; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_15; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_16; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_17; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_18; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_19; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_20; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_21; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_22; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_23; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_24; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_25; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_26; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_27; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_28; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_29; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_30; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_31; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_32; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_33; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_34; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_35; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_36; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_37; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_38; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_39; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_40; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_41; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_42; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_43; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_44; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_45; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_46; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_47; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_48; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_49; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_50; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_51; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_52; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_53; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_54; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_55; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_56; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_57; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_58; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_59; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_60; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_61; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_62; // @[BuildingBlockNew.scala 84:24]
  wire [3:0] ingress1_io_out64_63; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_0; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_1; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_2; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_3; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_4; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_5; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_6; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_7; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_8; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_9; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_10; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_11; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_12; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_13; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_14; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_15; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_16; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_17; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_18; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_19; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_20; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_21; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_22; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_23; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_24; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_25; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_26; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_27; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_28; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_29; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_30; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_31; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_32; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_33; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_34; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_35; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_36; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_37; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_38; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_39; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_40; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_41; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_42; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_43; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_44; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_45; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_46; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_47; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_48; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_49; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_50; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_51; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_52; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_53; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_54; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_55; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_56; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_57; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_58; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_59; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_60; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_61; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_62; // @[BuildingBlockNew.scala 84:24]
  wire  ingress1_io_validout64_63; // @[BuildingBlockNew.scala 84:24]
  wire [7:0] ingress1_io_addrout; // @[BuildingBlockNew.scala 84:24]
  wire [127:0] ingress1_io_ctrl; // @[BuildingBlockNew.scala 84:24]
  wire  ingress2_clock; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_0; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_1; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_2; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_3; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_4; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_5; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_6; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_7; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_8; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_9; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_10; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_11; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_12; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_13; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_14; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_15; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_16; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_17; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_18; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_19; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_20; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_21; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_22; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_23; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_24; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_25; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_26; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_27; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_28; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_29; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_30; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_31; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_32; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_33; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_34; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_35; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_36; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_37; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_38; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_39; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_40; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_41; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_42; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_43; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_44; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_45; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_46; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_47; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_48; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_49; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_50; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_51; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_52; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_53; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_54; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_55; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_56; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_57; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_58; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_59; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_60; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_61; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_62; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_in64_63; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_0; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_1; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_2; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_3; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_4; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_5; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_6; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_7; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_8; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_9; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_10; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_11; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_12; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_13; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_14; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_15; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_16; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_17; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_18; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_19; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_20; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_21; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_22; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_23; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_24; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_25; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_26; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_27; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_28; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_29; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_30; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_31; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_32; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_33; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_34; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_35; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_36; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_37; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_38; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_39; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_40; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_41; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_42; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_43; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_44; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_45; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_46; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_47; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_48; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_49; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_50; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_51; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_52; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_53; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_54; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_55; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_56; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_57; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_58; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_59; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_60; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_61; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_62; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validin64_63; // @[BuildingBlockNew.scala 85:24]
  wire [7:0] ingress2_io_addrin; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_0; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_1; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_2; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_3; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_4; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_5; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_6; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_7; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_8; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_9; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_10; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_11; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_12; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_13; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_14; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_15; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_16; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_17; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_18; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_19; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_20; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_21; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_22; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_23; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_24; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_25; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_26; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_27; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_28; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_29; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_30; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_31; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_32; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_33; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_34; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_35; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_36; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_37; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_38; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_39; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_40; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_41; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_42; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_43; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_44; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_45; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_46; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_47; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_48; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_49; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_50; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_51; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_52; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_53; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_54; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_55; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_56; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_57; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_58; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_59; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_60; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_61; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_62; // @[BuildingBlockNew.scala 85:24]
  wire [3:0] ingress2_io_out64_63; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_0; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_1; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_2; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_3; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_4; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_5; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_6; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_7; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_8; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_9; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_10; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_11; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_12; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_13; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_14; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_15; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_16; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_17; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_18; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_19; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_20; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_21; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_22; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_23; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_24; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_25; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_26; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_27; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_28; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_29; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_30; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_31; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_32; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_33; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_34; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_35; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_36; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_37; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_38; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_39; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_40; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_41; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_42; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_43; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_44; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_45; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_46; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_47; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_48; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_49; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_50; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_51; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_52; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_53; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_54; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_55; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_56; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_57; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_58; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_59; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_60; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_61; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_62; // @[BuildingBlockNew.scala 85:24]
  wire  ingress2_io_validout64_63; // @[BuildingBlockNew.scala 85:24]
  wire [7:0] ingress2_io_addrout; // @[BuildingBlockNew.scala 85:24]
  wire [127:0] ingress2_io_ctrl; // @[BuildingBlockNew.scala 85:24]
  wire  middle_clock; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_0; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_1; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_2; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_3; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_4; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_5; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_6; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_7; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_8; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_9; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_10; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_11; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_12; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_13; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_14; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_15; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_16; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_17; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_18; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_19; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_20; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_21; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_22; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_23; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_24; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_25; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_26; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_27; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_28; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_29; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_30; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_31; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_32; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_33; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_34; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_35; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_36; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_37; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_38; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_39; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_40; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_41; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_42; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_43; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_44; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_45; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_46; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_47; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_48; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_49; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_50; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_51; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_52; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_53; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_54; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_55; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_56; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_57; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_58; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_59; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_60; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_61; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_62; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_in64_63; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_0; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_1; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_2; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_3; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_4; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_5; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_6; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_7; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_8; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_9; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_10; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_11; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_12; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_13; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_14; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_15; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_16; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_17; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_18; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_19; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_20; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_21; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_22; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_23; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_24; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_25; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_26; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_27; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_28; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_29; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_30; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_31; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_32; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_33; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_34; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_35; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_36; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_37; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_38; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_39; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_40; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_41; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_42; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_43; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_44; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_45; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_46; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_47; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_48; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_49; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_50; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_51; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_52; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_53; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_54; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_55; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_56; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_57; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_58; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_59; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_60; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_61; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_62; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validin64_63; // @[BuildingBlockNew.scala 86:22]
  wire [7:0] middle_io_addrin; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_0; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_1; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_2; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_3; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_4; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_5; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_6; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_7; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_8; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_9; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_10; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_11; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_12; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_13; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_14; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_15; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_16; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_17; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_18; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_19; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_20; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_21; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_22; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_23; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_24; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_25; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_26; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_27; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_28; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_29; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_30; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_31; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_32; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_33; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_34; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_35; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_36; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_37; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_38; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_39; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_40; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_41; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_42; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_43; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_44; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_45; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_46; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_47; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_48; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_49; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_50; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_51; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_52; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_53; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_54; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_55; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_56; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_57; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_58; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_59; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_60; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_61; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_62; // @[BuildingBlockNew.scala 86:22]
  wire [3:0] middle_io_out64_63; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_0; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_1; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_2; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_3; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_4; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_5; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_6; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_7; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_8; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_9; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_10; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_11; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_12; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_13; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_14; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_15; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_16; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_17; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_18; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_19; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_20; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_21; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_22; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_23; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_24; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_25; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_26; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_27; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_28; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_29; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_30; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_31; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_32; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_33; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_34; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_35; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_36; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_37; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_38; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_39; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_40; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_41; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_42; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_43; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_44; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_45; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_46; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_47; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_48; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_49; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_50; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_51; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_52; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_53; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_54; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_55; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_56; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_57; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_58; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_59; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_60; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_61; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_62; // @[BuildingBlockNew.scala 86:22]
  wire  middle_io_validout64_63; // @[BuildingBlockNew.scala 86:22]
  wire [7:0] middle_io_addrout; // @[BuildingBlockNew.scala 86:22]
  wire [127:0] middle_io_ctrl; // @[BuildingBlockNew.scala 86:22]
  wire  egress1_clock; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_0; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_1; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_2; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_3; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_4; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_5; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_6; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_7; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_8; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_9; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_10; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_11; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_12; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_13; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_14; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_15; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_16; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_17; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_18; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_19; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_20; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_21; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_22; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_23; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_24; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_25; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_26; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_27; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_28; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_29; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_30; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_31; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_32; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_33; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_34; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_35; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_36; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_37; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_38; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_39; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_40; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_41; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_42; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_43; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_44; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_45; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_46; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_47; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_48; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_49; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_50; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_51; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_52; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_53; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_54; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_55; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_56; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_57; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_58; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_59; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_60; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_61; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_62; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_in64_63; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_0; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_1; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_2; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_3; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_4; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_5; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_6; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_7; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_8; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_9; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_10; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_11; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_12; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_13; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_14; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_15; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_16; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_17; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_18; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_19; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_20; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_21; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_22; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_23; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_24; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_25; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_26; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_27; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_28; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_29; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_30; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_31; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_32; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_33; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_34; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_35; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_36; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_37; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_38; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_39; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_40; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_41; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_42; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_43; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_44; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_45; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_46; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_47; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_48; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_49; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_50; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_51; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_52; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_53; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_54; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_55; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_56; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_57; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_58; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_59; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_60; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_61; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_62; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validin64_63; // @[BuildingBlockNew.scala 87:23]
  wire [7:0] egress1_io_addrin; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_0; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_1; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_2; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_3; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_4; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_5; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_6; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_7; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_8; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_9; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_10; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_11; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_12; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_13; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_14; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_15; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_16; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_17; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_18; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_19; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_20; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_21; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_22; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_23; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_24; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_25; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_26; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_27; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_28; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_29; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_30; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_31; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_32; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_33; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_34; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_35; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_36; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_37; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_38; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_39; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_40; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_41; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_42; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_43; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_44; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_45; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_46; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_47; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_48; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_49; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_50; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_51; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_52; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_53; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_54; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_55; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_56; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_57; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_58; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_59; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_60; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_61; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_62; // @[BuildingBlockNew.scala 87:23]
  wire [3:0] egress1_io_out64_63; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_0; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_1; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_2; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_3; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_4; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_5; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_6; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_7; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_8; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_9; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_10; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_11; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_12; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_13; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_14; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_15; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_16; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_17; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_18; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_19; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_20; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_21; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_22; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_23; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_24; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_25; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_26; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_27; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_28; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_29; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_30; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_31; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_32; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_33; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_34; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_35; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_36; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_37; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_38; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_39; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_40; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_41; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_42; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_43; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_44; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_45; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_46; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_47; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_48; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_49; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_50; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_51; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_52; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_53; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_54; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_55; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_56; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_57; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_58; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_59; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_60; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_61; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_62; // @[BuildingBlockNew.scala 87:23]
  wire  egress1_io_validout64_63; // @[BuildingBlockNew.scala 87:23]
  wire [7:0] egress1_io_addrout; // @[BuildingBlockNew.scala 87:23]
  wire [127:0] egress1_io_ctrl; // @[BuildingBlockNew.scala 87:23]
  wire  egress2_clock; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_0; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_1; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_2; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_3; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_4; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_5; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_6; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_7; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_8; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_9; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_10; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_11; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_12; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_13; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_14; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_15; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_16; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_17; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_18; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_19; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_20; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_21; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_22; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_23; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_24; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_25; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_26; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_27; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_28; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_29; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_30; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_31; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_32; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_33; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_34; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_35; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_36; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_37; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_38; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_39; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_40; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_41; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_42; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_43; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_44; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_45; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_46; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_47; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_48; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_49; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_50; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_51; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_52; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_53; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_54; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_55; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_56; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_57; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_58; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_59; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_60; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_61; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_62; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_in64_63; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_0; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_1; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_2; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_3; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_4; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_5; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_6; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_7; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_8; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_9; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_10; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_11; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_12; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_13; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_14; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_15; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_16; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_17; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_18; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_19; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_20; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_21; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_22; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_23; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_24; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_25; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_26; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_27; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_28; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_29; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_30; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_31; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_32; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_33; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_34; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_35; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_36; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_37; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_38; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_39; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_40; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_41; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_42; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_43; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_44; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_45; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_46; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_47; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_48; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_49; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_50; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_51; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_52; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_53; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_54; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_55; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_56; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_57; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_58; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_59; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_60; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_61; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_62; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validin64_63; // @[BuildingBlockNew.scala 88:23]
  wire [7:0] egress2_io_addrin; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_0; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_1; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_2; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_3; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_4; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_5; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_6; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_7; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_8; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_9; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_10; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_11; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_12; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_13; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_14; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_15; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_16; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_17; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_18; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_19; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_20; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_21; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_22; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_23; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_24; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_25; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_26; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_27; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_28; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_29; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_30; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_31; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_32; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_33; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_34; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_35; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_36; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_37; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_38; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_39; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_40; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_41; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_42; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_43; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_44; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_45; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_46; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_47; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_48; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_49; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_50; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_51; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_52; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_53; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_54; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_55; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_56; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_57; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_58; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_59; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_60; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_61; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_62; // @[BuildingBlockNew.scala 88:23]
  wire [3:0] egress2_io_out64_63; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_0; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_1; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_2; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_3; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_4; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_5; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_6; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_7; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_8; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_9; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_10; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_11; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_12; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_13; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_14; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_15; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_16; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_17; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_18; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_19; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_20; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_21; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_22; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_23; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_24; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_25; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_26; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_27; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_28; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_29; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_30; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_31; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_32; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_33; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_34; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_35; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_36; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_37; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_38; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_39; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_40; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_41; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_42; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_43; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_44; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_45; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_46; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_47; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_48; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_49; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_50; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_51; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_52; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_53; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_54; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_55; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_56; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_57; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_58; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_59; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_60; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_61; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_62; // @[BuildingBlockNew.scala 88:23]
  wire  egress2_io_validout64_63; // @[BuildingBlockNew.scala 88:23]
  wire [7:0] egress2_io_addrout; // @[BuildingBlockNew.scala 88:23]
  wire [127:0] egress2_io_ctrl; // @[BuildingBlockNew.scala 88:23]
  reg [7:0] PC1; // @[BuildingBlockNew.scala 39:20]
  reg [7:0] PC2; // @[BuildingBlockNew.scala 40:20]
  reg [7:0] PC3; // @[BuildingBlockNew.scala 41:20]
  reg [7:0] PC4; // @[BuildingBlockNew.scala 42:20]
  reg [7:0] PC5; // @[BuildingBlockNew.scala 43:20]
  reg [7:0] PC6; // @[BuildingBlockNew.scala 44:20]
  reg [7:0] wrAddr1; // @[BuildingBlockNew.scala 45:24]
  reg [7:0] wrAddr2; // @[BuildingBlockNew.scala 46:24]
  reg [7:0] wrAddr3; // @[BuildingBlockNew.scala 47:24]
  reg [7:0] wrAddr4; // @[BuildingBlockNew.scala 48:24]
  reg [7:0] wrAddr5; // @[BuildingBlockNew.scala 49:24]
  reg [7:0] wrAddr6; // @[BuildingBlockNew.scala 50:24]
  wire [7:0] _wrAddr1_T_1 = wrAddr1 + 8'h1; // @[BuildingBlockNew.scala 226:24]
  wire [7:0] _wrAddr2_T_1 = wrAddr2 + 8'h1; // @[BuildingBlockNew.scala 235:24]
  wire [7:0] _wrAddr3_T_1 = wrAddr3 + 8'h1; // @[BuildingBlockNew.scala 244:24]
  wire [7:0] _wrAddr4_T_1 = wrAddr4 + 8'h1; // @[BuildingBlockNew.scala 253:24]
  wire [7:0] _wrAddr5_T_1 = wrAddr5 + 8'h1; // @[BuildingBlockNew.scala 262:24]
  wire [7:0] _wrAddr6_T_1 = wrAddr6 + 8'h1; // @[BuildingBlockNew.scala 271:24]
  PEcol peCol ( // @[BuildingBlockNew.scala 83:21]
    .clock(peCol_clock),
    .reset(peCol_reset),
    .io_d_in_0_a(peCol_io_d_in_0_a),
    .io_d_in_0_valid_a(peCol_io_d_in_0_valid_a),
    .io_d_in_0_b(peCol_io_d_in_0_b),
    .io_d_in_0_valid_b(peCol_io_d_in_0_valid_b),
    .io_d_in_1_a(peCol_io_d_in_1_a),
    .io_d_in_1_valid_a(peCol_io_d_in_1_valid_a),
    .io_d_in_1_b(peCol_io_d_in_1_b),
    .io_d_in_1_valid_b(peCol_io_d_in_1_valid_b),
    .io_d_in_2_a(peCol_io_d_in_2_a),
    .io_d_in_2_valid_a(peCol_io_d_in_2_valid_a),
    .io_d_in_2_b(peCol_io_d_in_2_b),
    .io_d_in_2_valid_b(peCol_io_d_in_2_valid_b),
    .io_d_in_3_a(peCol_io_d_in_3_a),
    .io_d_in_3_valid_a(peCol_io_d_in_3_valid_a),
    .io_d_in_3_b(peCol_io_d_in_3_b),
    .io_d_in_3_valid_b(peCol_io_d_in_3_valid_b),
    .io_d_in_4_a(peCol_io_d_in_4_a),
    .io_d_in_4_valid_a(peCol_io_d_in_4_valid_a),
    .io_d_in_4_b(peCol_io_d_in_4_b),
    .io_d_in_4_valid_b(peCol_io_d_in_4_valid_b),
    .io_d_in_5_a(peCol_io_d_in_5_a),
    .io_d_in_5_valid_a(peCol_io_d_in_5_valid_a),
    .io_d_in_5_b(peCol_io_d_in_5_b),
    .io_d_in_5_valid_b(peCol_io_d_in_5_valid_b),
    .io_d_in_6_a(peCol_io_d_in_6_a),
    .io_d_in_6_valid_a(peCol_io_d_in_6_valid_a),
    .io_d_in_6_b(peCol_io_d_in_6_b),
    .io_d_in_6_valid_b(peCol_io_d_in_6_valid_b),
    .io_d_in_7_a(peCol_io_d_in_7_a),
    .io_d_in_7_valid_a(peCol_io_d_in_7_valid_a),
    .io_d_in_7_b(peCol_io_d_in_7_b),
    .io_d_in_7_valid_b(peCol_io_d_in_7_valid_b),
    .io_d_in_8_a(peCol_io_d_in_8_a),
    .io_d_in_8_valid_a(peCol_io_d_in_8_valid_a),
    .io_d_in_8_b(peCol_io_d_in_8_b),
    .io_d_in_8_valid_b(peCol_io_d_in_8_valid_b),
    .io_d_in_9_a(peCol_io_d_in_9_a),
    .io_d_in_9_valid_a(peCol_io_d_in_9_valid_a),
    .io_d_in_9_b(peCol_io_d_in_9_b),
    .io_d_in_9_valid_b(peCol_io_d_in_9_valid_b),
    .io_d_in_10_a(peCol_io_d_in_10_a),
    .io_d_in_10_valid_a(peCol_io_d_in_10_valid_a),
    .io_d_in_10_b(peCol_io_d_in_10_b),
    .io_d_in_10_valid_b(peCol_io_d_in_10_valid_b),
    .io_d_in_11_a(peCol_io_d_in_11_a),
    .io_d_in_11_valid_a(peCol_io_d_in_11_valid_a),
    .io_d_in_11_b(peCol_io_d_in_11_b),
    .io_d_in_11_valid_b(peCol_io_d_in_11_valid_b),
    .io_d_in_12_a(peCol_io_d_in_12_a),
    .io_d_in_12_valid_a(peCol_io_d_in_12_valid_a),
    .io_d_in_12_b(peCol_io_d_in_12_b),
    .io_d_in_12_valid_b(peCol_io_d_in_12_valid_b),
    .io_d_in_13_a(peCol_io_d_in_13_a),
    .io_d_in_13_valid_a(peCol_io_d_in_13_valid_a),
    .io_d_in_13_b(peCol_io_d_in_13_b),
    .io_d_in_13_valid_b(peCol_io_d_in_13_valid_b),
    .io_d_in_14_a(peCol_io_d_in_14_a),
    .io_d_in_14_valid_a(peCol_io_d_in_14_valid_a),
    .io_d_in_14_b(peCol_io_d_in_14_b),
    .io_d_in_14_valid_b(peCol_io_d_in_14_valid_b),
    .io_d_in_15_a(peCol_io_d_in_15_a),
    .io_d_in_15_valid_a(peCol_io_d_in_15_valid_a),
    .io_d_in_15_b(peCol_io_d_in_15_b),
    .io_d_in_15_valid_b(peCol_io_d_in_15_valid_b),
    .io_d_in_16_a(peCol_io_d_in_16_a),
    .io_d_in_16_valid_a(peCol_io_d_in_16_valid_a),
    .io_d_in_16_b(peCol_io_d_in_16_b),
    .io_d_in_16_valid_b(peCol_io_d_in_16_valid_b),
    .io_d_in_17_a(peCol_io_d_in_17_a),
    .io_d_in_17_valid_a(peCol_io_d_in_17_valid_a),
    .io_d_in_17_b(peCol_io_d_in_17_b),
    .io_d_in_17_valid_b(peCol_io_d_in_17_valid_b),
    .io_d_in_18_a(peCol_io_d_in_18_a),
    .io_d_in_18_valid_a(peCol_io_d_in_18_valid_a),
    .io_d_in_18_b(peCol_io_d_in_18_b),
    .io_d_in_18_valid_b(peCol_io_d_in_18_valid_b),
    .io_d_in_19_a(peCol_io_d_in_19_a),
    .io_d_in_19_valid_a(peCol_io_d_in_19_valid_a),
    .io_d_in_19_b(peCol_io_d_in_19_b),
    .io_d_in_19_valid_b(peCol_io_d_in_19_valid_b),
    .io_d_in_20_a(peCol_io_d_in_20_a),
    .io_d_in_20_valid_a(peCol_io_d_in_20_valid_a),
    .io_d_in_20_b(peCol_io_d_in_20_b),
    .io_d_in_20_valid_b(peCol_io_d_in_20_valid_b),
    .io_d_in_21_a(peCol_io_d_in_21_a),
    .io_d_in_21_valid_a(peCol_io_d_in_21_valid_a),
    .io_d_in_21_b(peCol_io_d_in_21_b),
    .io_d_in_21_valid_b(peCol_io_d_in_21_valid_b),
    .io_d_in_22_a(peCol_io_d_in_22_a),
    .io_d_in_22_valid_a(peCol_io_d_in_22_valid_a),
    .io_d_in_22_b(peCol_io_d_in_22_b),
    .io_d_in_22_valid_b(peCol_io_d_in_22_valid_b),
    .io_d_in_23_a(peCol_io_d_in_23_a),
    .io_d_in_23_valid_a(peCol_io_d_in_23_valid_a),
    .io_d_in_23_b(peCol_io_d_in_23_b),
    .io_d_in_23_valid_b(peCol_io_d_in_23_valid_b),
    .io_d_in_24_a(peCol_io_d_in_24_a),
    .io_d_in_24_valid_a(peCol_io_d_in_24_valid_a),
    .io_d_in_24_b(peCol_io_d_in_24_b),
    .io_d_in_24_valid_b(peCol_io_d_in_24_valid_b),
    .io_d_in_25_a(peCol_io_d_in_25_a),
    .io_d_in_25_valid_a(peCol_io_d_in_25_valid_a),
    .io_d_in_25_b(peCol_io_d_in_25_b),
    .io_d_in_25_valid_b(peCol_io_d_in_25_valid_b),
    .io_d_in_26_a(peCol_io_d_in_26_a),
    .io_d_in_26_valid_a(peCol_io_d_in_26_valid_a),
    .io_d_in_26_b(peCol_io_d_in_26_b),
    .io_d_in_26_valid_b(peCol_io_d_in_26_valid_b),
    .io_d_in_27_a(peCol_io_d_in_27_a),
    .io_d_in_27_valid_a(peCol_io_d_in_27_valid_a),
    .io_d_in_27_b(peCol_io_d_in_27_b),
    .io_d_in_27_valid_b(peCol_io_d_in_27_valid_b),
    .io_d_in_28_a(peCol_io_d_in_28_a),
    .io_d_in_28_valid_a(peCol_io_d_in_28_valid_a),
    .io_d_in_28_b(peCol_io_d_in_28_b),
    .io_d_in_28_valid_b(peCol_io_d_in_28_valid_b),
    .io_d_in_29_a(peCol_io_d_in_29_a),
    .io_d_in_29_valid_a(peCol_io_d_in_29_valid_a),
    .io_d_in_29_b(peCol_io_d_in_29_b),
    .io_d_in_29_valid_b(peCol_io_d_in_29_valid_b),
    .io_d_in_30_a(peCol_io_d_in_30_a),
    .io_d_in_30_valid_a(peCol_io_d_in_30_valid_a),
    .io_d_in_30_b(peCol_io_d_in_30_b),
    .io_d_in_30_valid_b(peCol_io_d_in_30_valid_b),
    .io_d_in_31_a(peCol_io_d_in_31_a),
    .io_d_in_31_valid_a(peCol_io_d_in_31_valid_a),
    .io_d_in_31_b(peCol_io_d_in_31_b),
    .io_d_in_31_valid_b(peCol_io_d_in_31_valid_b),
    .io_d_out_0_a(peCol_io_d_out_0_a),
    .io_d_out_0_valid_a(peCol_io_d_out_0_valid_a),
    .io_d_out_0_b(peCol_io_d_out_0_b),
    .io_d_out_0_valid_b(peCol_io_d_out_0_valid_b),
    .io_d_out_1_a(peCol_io_d_out_1_a),
    .io_d_out_1_valid_a(peCol_io_d_out_1_valid_a),
    .io_d_out_1_b(peCol_io_d_out_1_b),
    .io_d_out_1_valid_b(peCol_io_d_out_1_valid_b),
    .io_d_out_2_a(peCol_io_d_out_2_a),
    .io_d_out_2_valid_a(peCol_io_d_out_2_valid_a),
    .io_d_out_2_b(peCol_io_d_out_2_b),
    .io_d_out_2_valid_b(peCol_io_d_out_2_valid_b),
    .io_d_out_3_a(peCol_io_d_out_3_a),
    .io_d_out_3_valid_a(peCol_io_d_out_3_valid_a),
    .io_d_out_3_b(peCol_io_d_out_3_b),
    .io_d_out_3_valid_b(peCol_io_d_out_3_valid_b),
    .io_d_out_4_a(peCol_io_d_out_4_a),
    .io_d_out_4_valid_a(peCol_io_d_out_4_valid_a),
    .io_d_out_4_b(peCol_io_d_out_4_b),
    .io_d_out_4_valid_b(peCol_io_d_out_4_valid_b),
    .io_d_out_5_a(peCol_io_d_out_5_a),
    .io_d_out_5_valid_a(peCol_io_d_out_5_valid_a),
    .io_d_out_5_b(peCol_io_d_out_5_b),
    .io_d_out_5_valid_b(peCol_io_d_out_5_valid_b),
    .io_d_out_6_a(peCol_io_d_out_6_a),
    .io_d_out_6_valid_a(peCol_io_d_out_6_valid_a),
    .io_d_out_6_b(peCol_io_d_out_6_b),
    .io_d_out_6_valid_b(peCol_io_d_out_6_valid_b),
    .io_d_out_7_a(peCol_io_d_out_7_a),
    .io_d_out_7_valid_a(peCol_io_d_out_7_valid_a),
    .io_d_out_7_b(peCol_io_d_out_7_b),
    .io_d_out_7_valid_b(peCol_io_d_out_7_valid_b),
    .io_d_out_8_a(peCol_io_d_out_8_a),
    .io_d_out_8_valid_a(peCol_io_d_out_8_valid_a),
    .io_d_out_8_b(peCol_io_d_out_8_b),
    .io_d_out_8_valid_b(peCol_io_d_out_8_valid_b),
    .io_d_out_9_a(peCol_io_d_out_9_a),
    .io_d_out_9_valid_a(peCol_io_d_out_9_valid_a),
    .io_d_out_9_b(peCol_io_d_out_9_b),
    .io_d_out_9_valid_b(peCol_io_d_out_9_valid_b),
    .io_d_out_10_a(peCol_io_d_out_10_a),
    .io_d_out_10_valid_a(peCol_io_d_out_10_valid_a),
    .io_d_out_10_b(peCol_io_d_out_10_b),
    .io_d_out_10_valid_b(peCol_io_d_out_10_valid_b),
    .io_d_out_11_a(peCol_io_d_out_11_a),
    .io_d_out_11_valid_a(peCol_io_d_out_11_valid_a),
    .io_d_out_11_b(peCol_io_d_out_11_b),
    .io_d_out_11_valid_b(peCol_io_d_out_11_valid_b),
    .io_d_out_12_a(peCol_io_d_out_12_a),
    .io_d_out_12_valid_a(peCol_io_d_out_12_valid_a),
    .io_d_out_12_b(peCol_io_d_out_12_b),
    .io_d_out_12_valid_b(peCol_io_d_out_12_valid_b),
    .io_d_out_13_a(peCol_io_d_out_13_a),
    .io_d_out_13_valid_a(peCol_io_d_out_13_valid_a),
    .io_d_out_13_b(peCol_io_d_out_13_b),
    .io_d_out_13_valid_b(peCol_io_d_out_13_valid_b),
    .io_d_out_14_a(peCol_io_d_out_14_a),
    .io_d_out_14_valid_a(peCol_io_d_out_14_valid_a),
    .io_d_out_14_b(peCol_io_d_out_14_b),
    .io_d_out_14_valid_b(peCol_io_d_out_14_valid_b),
    .io_d_out_15_a(peCol_io_d_out_15_a),
    .io_d_out_15_valid_a(peCol_io_d_out_15_valid_a),
    .io_d_out_15_b(peCol_io_d_out_15_b),
    .io_d_out_15_valid_b(peCol_io_d_out_15_valid_b),
    .io_d_out_16_a(peCol_io_d_out_16_a),
    .io_d_out_16_valid_a(peCol_io_d_out_16_valid_a),
    .io_d_out_16_b(peCol_io_d_out_16_b),
    .io_d_out_16_valid_b(peCol_io_d_out_16_valid_b),
    .io_d_out_17_a(peCol_io_d_out_17_a),
    .io_d_out_17_valid_a(peCol_io_d_out_17_valid_a),
    .io_d_out_17_b(peCol_io_d_out_17_b),
    .io_d_out_17_valid_b(peCol_io_d_out_17_valid_b),
    .io_d_out_18_a(peCol_io_d_out_18_a),
    .io_d_out_18_valid_a(peCol_io_d_out_18_valid_a),
    .io_d_out_18_b(peCol_io_d_out_18_b),
    .io_d_out_18_valid_b(peCol_io_d_out_18_valid_b),
    .io_d_out_19_a(peCol_io_d_out_19_a),
    .io_d_out_19_valid_a(peCol_io_d_out_19_valid_a),
    .io_d_out_19_b(peCol_io_d_out_19_b),
    .io_d_out_19_valid_b(peCol_io_d_out_19_valid_b),
    .io_d_out_20_a(peCol_io_d_out_20_a),
    .io_d_out_20_valid_a(peCol_io_d_out_20_valid_a),
    .io_d_out_20_b(peCol_io_d_out_20_b),
    .io_d_out_20_valid_b(peCol_io_d_out_20_valid_b),
    .io_d_out_21_a(peCol_io_d_out_21_a),
    .io_d_out_21_valid_a(peCol_io_d_out_21_valid_a),
    .io_d_out_21_b(peCol_io_d_out_21_b),
    .io_d_out_21_valid_b(peCol_io_d_out_21_valid_b),
    .io_d_out_22_a(peCol_io_d_out_22_a),
    .io_d_out_22_valid_a(peCol_io_d_out_22_valid_a),
    .io_d_out_22_b(peCol_io_d_out_22_b),
    .io_d_out_22_valid_b(peCol_io_d_out_22_valid_b),
    .io_d_out_23_a(peCol_io_d_out_23_a),
    .io_d_out_23_valid_a(peCol_io_d_out_23_valid_a),
    .io_d_out_23_b(peCol_io_d_out_23_b),
    .io_d_out_23_valid_b(peCol_io_d_out_23_valid_b),
    .io_d_out_24_a(peCol_io_d_out_24_a),
    .io_d_out_24_valid_a(peCol_io_d_out_24_valid_a),
    .io_d_out_24_b(peCol_io_d_out_24_b),
    .io_d_out_24_valid_b(peCol_io_d_out_24_valid_b),
    .io_d_out_25_a(peCol_io_d_out_25_a),
    .io_d_out_25_valid_a(peCol_io_d_out_25_valid_a),
    .io_d_out_25_b(peCol_io_d_out_25_b),
    .io_d_out_25_valid_b(peCol_io_d_out_25_valid_b),
    .io_d_out_26_a(peCol_io_d_out_26_a),
    .io_d_out_26_valid_a(peCol_io_d_out_26_valid_a),
    .io_d_out_26_b(peCol_io_d_out_26_b),
    .io_d_out_26_valid_b(peCol_io_d_out_26_valid_b),
    .io_d_out_27_a(peCol_io_d_out_27_a),
    .io_d_out_27_valid_a(peCol_io_d_out_27_valid_a),
    .io_d_out_27_b(peCol_io_d_out_27_b),
    .io_d_out_27_valid_b(peCol_io_d_out_27_valid_b),
    .io_d_out_28_a(peCol_io_d_out_28_a),
    .io_d_out_28_valid_a(peCol_io_d_out_28_valid_a),
    .io_d_out_28_b(peCol_io_d_out_28_b),
    .io_d_out_28_valid_b(peCol_io_d_out_28_valid_b),
    .io_d_out_29_a(peCol_io_d_out_29_a),
    .io_d_out_29_valid_a(peCol_io_d_out_29_valid_a),
    .io_d_out_29_b(peCol_io_d_out_29_b),
    .io_d_out_29_valid_b(peCol_io_d_out_29_valid_b),
    .io_d_out_30_a(peCol_io_d_out_30_a),
    .io_d_out_30_valid_a(peCol_io_d_out_30_valid_a),
    .io_d_out_30_b(peCol_io_d_out_30_b),
    .io_d_out_30_valid_b(peCol_io_d_out_30_valid_b),
    .io_d_out_31_a(peCol_io_d_out_31_a),
    .io_d_out_31_valid_a(peCol_io_d_out_31_valid_a),
    .io_d_out_31_b(peCol_io_d_out_31_b),
    .io_d_out_31_valid_b(peCol_io_d_out_31_valid_b),
    .io_addrin(peCol_io_addrin),
    .io_addrout(peCol_io_addrout),
    .io_instr(peCol_io_instr)
  );
  CLOSingress1 ingress1 ( // @[BuildingBlockNew.scala 84:24]
    .clock(ingress1_clock),
    .io_in64_0(ingress1_io_in64_0),
    .io_in64_1(ingress1_io_in64_1),
    .io_in64_2(ingress1_io_in64_2),
    .io_in64_3(ingress1_io_in64_3),
    .io_in64_4(ingress1_io_in64_4),
    .io_in64_5(ingress1_io_in64_5),
    .io_in64_6(ingress1_io_in64_6),
    .io_in64_7(ingress1_io_in64_7),
    .io_in64_8(ingress1_io_in64_8),
    .io_in64_9(ingress1_io_in64_9),
    .io_in64_10(ingress1_io_in64_10),
    .io_in64_11(ingress1_io_in64_11),
    .io_in64_12(ingress1_io_in64_12),
    .io_in64_13(ingress1_io_in64_13),
    .io_in64_14(ingress1_io_in64_14),
    .io_in64_15(ingress1_io_in64_15),
    .io_in64_16(ingress1_io_in64_16),
    .io_in64_17(ingress1_io_in64_17),
    .io_in64_18(ingress1_io_in64_18),
    .io_in64_19(ingress1_io_in64_19),
    .io_in64_20(ingress1_io_in64_20),
    .io_in64_21(ingress1_io_in64_21),
    .io_in64_22(ingress1_io_in64_22),
    .io_in64_23(ingress1_io_in64_23),
    .io_in64_24(ingress1_io_in64_24),
    .io_in64_25(ingress1_io_in64_25),
    .io_in64_26(ingress1_io_in64_26),
    .io_in64_27(ingress1_io_in64_27),
    .io_in64_28(ingress1_io_in64_28),
    .io_in64_29(ingress1_io_in64_29),
    .io_in64_30(ingress1_io_in64_30),
    .io_in64_31(ingress1_io_in64_31),
    .io_in64_32(ingress1_io_in64_32),
    .io_in64_33(ingress1_io_in64_33),
    .io_in64_34(ingress1_io_in64_34),
    .io_in64_35(ingress1_io_in64_35),
    .io_in64_36(ingress1_io_in64_36),
    .io_in64_37(ingress1_io_in64_37),
    .io_in64_38(ingress1_io_in64_38),
    .io_in64_39(ingress1_io_in64_39),
    .io_in64_40(ingress1_io_in64_40),
    .io_in64_41(ingress1_io_in64_41),
    .io_in64_42(ingress1_io_in64_42),
    .io_in64_43(ingress1_io_in64_43),
    .io_in64_44(ingress1_io_in64_44),
    .io_in64_45(ingress1_io_in64_45),
    .io_in64_46(ingress1_io_in64_46),
    .io_in64_47(ingress1_io_in64_47),
    .io_in64_48(ingress1_io_in64_48),
    .io_in64_49(ingress1_io_in64_49),
    .io_in64_50(ingress1_io_in64_50),
    .io_in64_51(ingress1_io_in64_51),
    .io_in64_52(ingress1_io_in64_52),
    .io_in64_53(ingress1_io_in64_53),
    .io_in64_54(ingress1_io_in64_54),
    .io_in64_55(ingress1_io_in64_55),
    .io_in64_56(ingress1_io_in64_56),
    .io_in64_57(ingress1_io_in64_57),
    .io_in64_58(ingress1_io_in64_58),
    .io_in64_59(ingress1_io_in64_59),
    .io_in64_60(ingress1_io_in64_60),
    .io_in64_61(ingress1_io_in64_61),
    .io_in64_62(ingress1_io_in64_62),
    .io_in64_63(ingress1_io_in64_63),
    .io_validin64_0(ingress1_io_validin64_0),
    .io_validin64_1(ingress1_io_validin64_1),
    .io_validin64_2(ingress1_io_validin64_2),
    .io_validin64_3(ingress1_io_validin64_3),
    .io_validin64_4(ingress1_io_validin64_4),
    .io_validin64_5(ingress1_io_validin64_5),
    .io_validin64_6(ingress1_io_validin64_6),
    .io_validin64_7(ingress1_io_validin64_7),
    .io_validin64_8(ingress1_io_validin64_8),
    .io_validin64_9(ingress1_io_validin64_9),
    .io_validin64_10(ingress1_io_validin64_10),
    .io_validin64_11(ingress1_io_validin64_11),
    .io_validin64_12(ingress1_io_validin64_12),
    .io_validin64_13(ingress1_io_validin64_13),
    .io_validin64_14(ingress1_io_validin64_14),
    .io_validin64_15(ingress1_io_validin64_15),
    .io_validin64_16(ingress1_io_validin64_16),
    .io_validin64_17(ingress1_io_validin64_17),
    .io_validin64_18(ingress1_io_validin64_18),
    .io_validin64_19(ingress1_io_validin64_19),
    .io_validin64_20(ingress1_io_validin64_20),
    .io_validin64_21(ingress1_io_validin64_21),
    .io_validin64_22(ingress1_io_validin64_22),
    .io_validin64_23(ingress1_io_validin64_23),
    .io_validin64_24(ingress1_io_validin64_24),
    .io_validin64_25(ingress1_io_validin64_25),
    .io_validin64_26(ingress1_io_validin64_26),
    .io_validin64_27(ingress1_io_validin64_27),
    .io_validin64_28(ingress1_io_validin64_28),
    .io_validin64_29(ingress1_io_validin64_29),
    .io_validin64_30(ingress1_io_validin64_30),
    .io_validin64_31(ingress1_io_validin64_31),
    .io_validin64_32(ingress1_io_validin64_32),
    .io_validin64_33(ingress1_io_validin64_33),
    .io_validin64_34(ingress1_io_validin64_34),
    .io_validin64_35(ingress1_io_validin64_35),
    .io_validin64_36(ingress1_io_validin64_36),
    .io_validin64_37(ingress1_io_validin64_37),
    .io_validin64_38(ingress1_io_validin64_38),
    .io_validin64_39(ingress1_io_validin64_39),
    .io_validin64_40(ingress1_io_validin64_40),
    .io_validin64_41(ingress1_io_validin64_41),
    .io_validin64_42(ingress1_io_validin64_42),
    .io_validin64_43(ingress1_io_validin64_43),
    .io_validin64_44(ingress1_io_validin64_44),
    .io_validin64_45(ingress1_io_validin64_45),
    .io_validin64_46(ingress1_io_validin64_46),
    .io_validin64_47(ingress1_io_validin64_47),
    .io_validin64_48(ingress1_io_validin64_48),
    .io_validin64_49(ingress1_io_validin64_49),
    .io_validin64_50(ingress1_io_validin64_50),
    .io_validin64_51(ingress1_io_validin64_51),
    .io_validin64_52(ingress1_io_validin64_52),
    .io_validin64_53(ingress1_io_validin64_53),
    .io_validin64_54(ingress1_io_validin64_54),
    .io_validin64_55(ingress1_io_validin64_55),
    .io_validin64_56(ingress1_io_validin64_56),
    .io_validin64_57(ingress1_io_validin64_57),
    .io_validin64_58(ingress1_io_validin64_58),
    .io_validin64_59(ingress1_io_validin64_59),
    .io_validin64_60(ingress1_io_validin64_60),
    .io_validin64_61(ingress1_io_validin64_61),
    .io_validin64_62(ingress1_io_validin64_62),
    .io_validin64_63(ingress1_io_validin64_63),
    .io_addrin(ingress1_io_addrin),
    .io_out64_0(ingress1_io_out64_0),
    .io_out64_1(ingress1_io_out64_1),
    .io_out64_2(ingress1_io_out64_2),
    .io_out64_3(ingress1_io_out64_3),
    .io_out64_4(ingress1_io_out64_4),
    .io_out64_5(ingress1_io_out64_5),
    .io_out64_6(ingress1_io_out64_6),
    .io_out64_7(ingress1_io_out64_7),
    .io_out64_8(ingress1_io_out64_8),
    .io_out64_9(ingress1_io_out64_9),
    .io_out64_10(ingress1_io_out64_10),
    .io_out64_11(ingress1_io_out64_11),
    .io_out64_12(ingress1_io_out64_12),
    .io_out64_13(ingress1_io_out64_13),
    .io_out64_14(ingress1_io_out64_14),
    .io_out64_15(ingress1_io_out64_15),
    .io_out64_16(ingress1_io_out64_16),
    .io_out64_17(ingress1_io_out64_17),
    .io_out64_18(ingress1_io_out64_18),
    .io_out64_19(ingress1_io_out64_19),
    .io_out64_20(ingress1_io_out64_20),
    .io_out64_21(ingress1_io_out64_21),
    .io_out64_22(ingress1_io_out64_22),
    .io_out64_23(ingress1_io_out64_23),
    .io_out64_24(ingress1_io_out64_24),
    .io_out64_25(ingress1_io_out64_25),
    .io_out64_26(ingress1_io_out64_26),
    .io_out64_27(ingress1_io_out64_27),
    .io_out64_28(ingress1_io_out64_28),
    .io_out64_29(ingress1_io_out64_29),
    .io_out64_30(ingress1_io_out64_30),
    .io_out64_31(ingress1_io_out64_31),
    .io_out64_32(ingress1_io_out64_32),
    .io_out64_33(ingress1_io_out64_33),
    .io_out64_34(ingress1_io_out64_34),
    .io_out64_35(ingress1_io_out64_35),
    .io_out64_36(ingress1_io_out64_36),
    .io_out64_37(ingress1_io_out64_37),
    .io_out64_38(ingress1_io_out64_38),
    .io_out64_39(ingress1_io_out64_39),
    .io_out64_40(ingress1_io_out64_40),
    .io_out64_41(ingress1_io_out64_41),
    .io_out64_42(ingress1_io_out64_42),
    .io_out64_43(ingress1_io_out64_43),
    .io_out64_44(ingress1_io_out64_44),
    .io_out64_45(ingress1_io_out64_45),
    .io_out64_46(ingress1_io_out64_46),
    .io_out64_47(ingress1_io_out64_47),
    .io_out64_48(ingress1_io_out64_48),
    .io_out64_49(ingress1_io_out64_49),
    .io_out64_50(ingress1_io_out64_50),
    .io_out64_51(ingress1_io_out64_51),
    .io_out64_52(ingress1_io_out64_52),
    .io_out64_53(ingress1_io_out64_53),
    .io_out64_54(ingress1_io_out64_54),
    .io_out64_55(ingress1_io_out64_55),
    .io_out64_56(ingress1_io_out64_56),
    .io_out64_57(ingress1_io_out64_57),
    .io_out64_58(ingress1_io_out64_58),
    .io_out64_59(ingress1_io_out64_59),
    .io_out64_60(ingress1_io_out64_60),
    .io_out64_61(ingress1_io_out64_61),
    .io_out64_62(ingress1_io_out64_62),
    .io_out64_63(ingress1_io_out64_63),
    .io_validout64_0(ingress1_io_validout64_0),
    .io_validout64_1(ingress1_io_validout64_1),
    .io_validout64_2(ingress1_io_validout64_2),
    .io_validout64_3(ingress1_io_validout64_3),
    .io_validout64_4(ingress1_io_validout64_4),
    .io_validout64_5(ingress1_io_validout64_5),
    .io_validout64_6(ingress1_io_validout64_6),
    .io_validout64_7(ingress1_io_validout64_7),
    .io_validout64_8(ingress1_io_validout64_8),
    .io_validout64_9(ingress1_io_validout64_9),
    .io_validout64_10(ingress1_io_validout64_10),
    .io_validout64_11(ingress1_io_validout64_11),
    .io_validout64_12(ingress1_io_validout64_12),
    .io_validout64_13(ingress1_io_validout64_13),
    .io_validout64_14(ingress1_io_validout64_14),
    .io_validout64_15(ingress1_io_validout64_15),
    .io_validout64_16(ingress1_io_validout64_16),
    .io_validout64_17(ingress1_io_validout64_17),
    .io_validout64_18(ingress1_io_validout64_18),
    .io_validout64_19(ingress1_io_validout64_19),
    .io_validout64_20(ingress1_io_validout64_20),
    .io_validout64_21(ingress1_io_validout64_21),
    .io_validout64_22(ingress1_io_validout64_22),
    .io_validout64_23(ingress1_io_validout64_23),
    .io_validout64_24(ingress1_io_validout64_24),
    .io_validout64_25(ingress1_io_validout64_25),
    .io_validout64_26(ingress1_io_validout64_26),
    .io_validout64_27(ingress1_io_validout64_27),
    .io_validout64_28(ingress1_io_validout64_28),
    .io_validout64_29(ingress1_io_validout64_29),
    .io_validout64_30(ingress1_io_validout64_30),
    .io_validout64_31(ingress1_io_validout64_31),
    .io_validout64_32(ingress1_io_validout64_32),
    .io_validout64_33(ingress1_io_validout64_33),
    .io_validout64_34(ingress1_io_validout64_34),
    .io_validout64_35(ingress1_io_validout64_35),
    .io_validout64_36(ingress1_io_validout64_36),
    .io_validout64_37(ingress1_io_validout64_37),
    .io_validout64_38(ingress1_io_validout64_38),
    .io_validout64_39(ingress1_io_validout64_39),
    .io_validout64_40(ingress1_io_validout64_40),
    .io_validout64_41(ingress1_io_validout64_41),
    .io_validout64_42(ingress1_io_validout64_42),
    .io_validout64_43(ingress1_io_validout64_43),
    .io_validout64_44(ingress1_io_validout64_44),
    .io_validout64_45(ingress1_io_validout64_45),
    .io_validout64_46(ingress1_io_validout64_46),
    .io_validout64_47(ingress1_io_validout64_47),
    .io_validout64_48(ingress1_io_validout64_48),
    .io_validout64_49(ingress1_io_validout64_49),
    .io_validout64_50(ingress1_io_validout64_50),
    .io_validout64_51(ingress1_io_validout64_51),
    .io_validout64_52(ingress1_io_validout64_52),
    .io_validout64_53(ingress1_io_validout64_53),
    .io_validout64_54(ingress1_io_validout64_54),
    .io_validout64_55(ingress1_io_validout64_55),
    .io_validout64_56(ingress1_io_validout64_56),
    .io_validout64_57(ingress1_io_validout64_57),
    .io_validout64_58(ingress1_io_validout64_58),
    .io_validout64_59(ingress1_io_validout64_59),
    .io_validout64_60(ingress1_io_validout64_60),
    .io_validout64_61(ingress1_io_validout64_61),
    .io_validout64_62(ingress1_io_validout64_62),
    .io_validout64_63(ingress1_io_validout64_63),
    .io_addrout(ingress1_io_addrout),
    .io_ctrl(ingress1_io_ctrl)
  );
  CLOSingress2 ingress2 ( // @[BuildingBlockNew.scala 85:24]
    .clock(ingress2_clock),
    .io_in64_0(ingress2_io_in64_0),
    .io_in64_1(ingress2_io_in64_1),
    .io_in64_2(ingress2_io_in64_2),
    .io_in64_3(ingress2_io_in64_3),
    .io_in64_4(ingress2_io_in64_4),
    .io_in64_5(ingress2_io_in64_5),
    .io_in64_6(ingress2_io_in64_6),
    .io_in64_7(ingress2_io_in64_7),
    .io_in64_8(ingress2_io_in64_8),
    .io_in64_9(ingress2_io_in64_9),
    .io_in64_10(ingress2_io_in64_10),
    .io_in64_11(ingress2_io_in64_11),
    .io_in64_12(ingress2_io_in64_12),
    .io_in64_13(ingress2_io_in64_13),
    .io_in64_14(ingress2_io_in64_14),
    .io_in64_15(ingress2_io_in64_15),
    .io_in64_16(ingress2_io_in64_16),
    .io_in64_17(ingress2_io_in64_17),
    .io_in64_18(ingress2_io_in64_18),
    .io_in64_19(ingress2_io_in64_19),
    .io_in64_20(ingress2_io_in64_20),
    .io_in64_21(ingress2_io_in64_21),
    .io_in64_22(ingress2_io_in64_22),
    .io_in64_23(ingress2_io_in64_23),
    .io_in64_24(ingress2_io_in64_24),
    .io_in64_25(ingress2_io_in64_25),
    .io_in64_26(ingress2_io_in64_26),
    .io_in64_27(ingress2_io_in64_27),
    .io_in64_28(ingress2_io_in64_28),
    .io_in64_29(ingress2_io_in64_29),
    .io_in64_30(ingress2_io_in64_30),
    .io_in64_31(ingress2_io_in64_31),
    .io_in64_32(ingress2_io_in64_32),
    .io_in64_33(ingress2_io_in64_33),
    .io_in64_34(ingress2_io_in64_34),
    .io_in64_35(ingress2_io_in64_35),
    .io_in64_36(ingress2_io_in64_36),
    .io_in64_37(ingress2_io_in64_37),
    .io_in64_38(ingress2_io_in64_38),
    .io_in64_39(ingress2_io_in64_39),
    .io_in64_40(ingress2_io_in64_40),
    .io_in64_41(ingress2_io_in64_41),
    .io_in64_42(ingress2_io_in64_42),
    .io_in64_43(ingress2_io_in64_43),
    .io_in64_44(ingress2_io_in64_44),
    .io_in64_45(ingress2_io_in64_45),
    .io_in64_46(ingress2_io_in64_46),
    .io_in64_47(ingress2_io_in64_47),
    .io_in64_48(ingress2_io_in64_48),
    .io_in64_49(ingress2_io_in64_49),
    .io_in64_50(ingress2_io_in64_50),
    .io_in64_51(ingress2_io_in64_51),
    .io_in64_52(ingress2_io_in64_52),
    .io_in64_53(ingress2_io_in64_53),
    .io_in64_54(ingress2_io_in64_54),
    .io_in64_55(ingress2_io_in64_55),
    .io_in64_56(ingress2_io_in64_56),
    .io_in64_57(ingress2_io_in64_57),
    .io_in64_58(ingress2_io_in64_58),
    .io_in64_59(ingress2_io_in64_59),
    .io_in64_60(ingress2_io_in64_60),
    .io_in64_61(ingress2_io_in64_61),
    .io_in64_62(ingress2_io_in64_62),
    .io_in64_63(ingress2_io_in64_63),
    .io_validin64_0(ingress2_io_validin64_0),
    .io_validin64_1(ingress2_io_validin64_1),
    .io_validin64_2(ingress2_io_validin64_2),
    .io_validin64_3(ingress2_io_validin64_3),
    .io_validin64_4(ingress2_io_validin64_4),
    .io_validin64_5(ingress2_io_validin64_5),
    .io_validin64_6(ingress2_io_validin64_6),
    .io_validin64_7(ingress2_io_validin64_7),
    .io_validin64_8(ingress2_io_validin64_8),
    .io_validin64_9(ingress2_io_validin64_9),
    .io_validin64_10(ingress2_io_validin64_10),
    .io_validin64_11(ingress2_io_validin64_11),
    .io_validin64_12(ingress2_io_validin64_12),
    .io_validin64_13(ingress2_io_validin64_13),
    .io_validin64_14(ingress2_io_validin64_14),
    .io_validin64_15(ingress2_io_validin64_15),
    .io_validin64_16(ingress2_io_validin64_16),
    .io_validin64_17(ingress2_io_validin64_17),
    .io_validin64_18(ingress2_io_validin64_18),
    .io_validin64_19(ingress2_io_validin64_19),
    .io_validin64_20(ingress2_io_validin64_20),
    .io_validin64_21(ingress2_io_validin64_21),
    .io_validin64_22(ingress2_io_validin64_22),
    .io_validin64_23(ingress2_io_validin64_23),
    .io_validin64_24(ingress2_io_validin64_24),
    .io_validin64_25(ingress2_io_validin64_25),
    .io_validin64_26(ingress2_io_validin64_26),
    .io_validin64_27(ingress2_io_validin64_27),
    .io_validin64_28(ingress2_io_validin64_28),
    .io_validin64_29(ingress2_io_validin64_29),
    .io_validin64_30(ingress2_io_validin64_30),
    .io_validin64_31(ingress2_io_validin64_31),
    .io_validin64_32(ingress2_io_validin64_32),
    .io_validin64_33(ingress2_io_validin64_33),
    .io_validin64_34(ingress2_io_validin64_34),
    .io_validin64_35(ingress2_io_validin64_35),
    .io_validin64_36(ingress2_io_validin64_36),
    .io_validin64_37(ingress2_io_validin64_37),
    .io_validin64_38(ingress2_io_validin64_38),
    .io_validin64_39(ingress2_io_validin64_39),
    .io_validin64_40(ingress2_io_validin64_40),
    .io_validin64_41(ingress2_io_validin64_41),
    .io_validin64_42(ingress2_io_validin64_42),
    .io_validin64_43(ingress2_io_validin64_43),
    .io_validin64_44(ingress2_io_validin64_44),
    .io_validin64_45(ingress2_io_validin64_45),
    .io_validin64_46(ingress2_io_validin64_46),
    .io_validin64_47(ingress2_io_validin64_47),
    .io_validin64_48(ingress2_io_validin64_48),
    .io_validin64_49(ingress2_io_validin64_49),
    .io_validin64_50(ingress2_io_validin64_50),
    .io_validin64_51(ingress2_io_validin64_51),
    .io_validin64_52(ingress2_io_validin64_52),
    .io_validin64_53(ingress2_io_validin64_53),
    .io_validin64_54(ingress2_io_validin64_54),
    .io_validin64_55(ingress2_io_validin64_55),
    .io_validin64_56(ingress2_io_validin64_56),
    .io_validin64_57(ingress2_io_validin64_57),
    .io_validin64_58(ingress2_io_validin64_58),
    .io_validin64_59(ingress2_io_validin64_59),
    .io_validin64_60(ingress2_io_validin64_60),
    .io_validin64_61(ingress2_io_validin64_61),
    .io_validin64_62(ingress2_io_validin64_62),
    .io_validin64_63(ingress2_io_validin64_63),
    .io_addrin(ingress2_io_addrin),
    .io_out64_0(ingress2_io_out64_0),
    .io_out64_1(ingress2_io_out64_1),
    .io_out64_2(ingress2_io_out64_2),
    .io_out64_3(ingress2_io_out64_3),
    .io_out64_4(ingress2_io_out64_4),
    .io_out64_5(ingress2_io_out64_5),
    .io_out64_6(ingress2_io_out64_6),
    .io_out64_7(ingress2_io_out64_7),
    .io_out64_8(ingress2_io_out64_8),
    .io_out64_9(ingress2_io_out64_9),
    .io_out64_10(ingress2_io_out64_10),
    .io_out64_11(ingress2_io_out64_11),
    .io_out64_12(ingress2_io_out64_12),
    .io_out64_13(ingress2_io_out64_13),
    .io_out64_14(ingress2_io_out64_14),
    .io_out64_15(ingress2_io_out64_15),
    .io_out64_16(ingress2_io_out64_16),
    .io_out64_17(ingress2_io_out64_17),
    .io_out64_18(ingress2_io_out64_18),
    .io_out64_19(ingress2_io_out64_19),
    .io_out64_20(ingress2_io_out64_20),
    .io_out64_21(ingress2_io_out64_21),
    .io_out64_22(ingress2_io_out64_22),
    .io_out64_23(ingress2_io_out64_23),
    .io_out64_24(ingress2_io_out64_24),
    .io_out64_25(ingress2_io_out64_25),
    .io_out64_26(ingress2_io_out64_26),
    .io_out64_27(ingress2_io_out64_27),
    .io_out64_28(ingress2_io_out64_28),
    .io_out64_29(ingress2_io_out64_29),
    .io_out64_30(ingress2_io_out64_30),
    .io_out64_31(ingress2_io_out64_31),
    .io_out64_32(ingress2_io_out64_32),
    .io_out64_33(ingress2_io_out64_33),
    .io_out64_34(ingress2_io_out64_34),
    .io_out64_35(ingress2_io_out64_35),
    .io_out64_36(ingress2_io_out64_36),
    .io_out64_37(ingress2_io_out64_37),
    .io_out64_38(ingress2_io_out64_38),
    .io_out64_39(ingress2_io_out64_39),
    .io_out64_40(ingress2_io_out64_40),
    .io_out64_41(ingress2_io_out64_41),
    .io_out64_42(ingress2_io_out64_42),
    .io_out64_43(ingress2_io_out64_43),
    .io_out64_44(ingress2_io_out64_44),
    .io_out64_45(ingress2_io_out64_45),
    .io_out64_46(ingress2_io_out64_46),
    .io_out64_47(ingress2_io_out64_47),
    .io_out64_48(ingress2_io_out64_48),
    .io_out64_49(ingress2_io_out64_49),
    .io_out64_50(ingress2_io_out64_50),
    .io_out64_51(ingress2_io_out64_51),
    .io_out64_52(ingress2_io_out64_52),
    .io_out64_53(ingress2_io_out64_53),
    .io_out64_54(ingress2_io_out64_54),
    .io_out64_55(ingress2_io_out64_55),
    .io_out64_56(ingress2_io_out64_56),
    .io_out64_57(ingress2_io_out64_57),
    .io_out64_58(ingress2_io_out64_58),
    .io_out64_59(ingress2_io_out64_59),
    .io_out64_60(ingress2_io_out64_60),
    .io_out64_61(ingress2_io_out64_61),
    .io_out64_62(ingress2_io_out64_62),
    .io_out64_63(ingress2_io_out64_63),
    .io_validout64_0(ingress2_io_validout64_0),
    .io_validout64_1(ingress2_io_validout64_1),
    .io_validout64_2(ingress2_io_validout64_2),
    .io_validout64_3(ingress2_io_validout64_3),
    .io_validout64_4(ingress2_io_validout64_4),
    .io_validout64_5(ingress2_io_validout64_5),
    .io_validout64_6(ingress2_io_validout64_6),
    .io_validout64_7(ingress2_io_validout64_7),
    .io_validout64_8(ingress2_io_validout64_8),
    .io_validout64_9(ingress2_io_validout64_9),
    .io_validout64_10(ingress2_io_validout64_10),
    .io_validout64_11(ingress2_io_validout64_11),
    .io_validout64_12(ingress2_io_validout64_12),
    .io_validout64_13(ingress2_io_validout64_13),
    .io_validout64_14(ingress2_io_validout64_14),
    .io_validout64_15(ingress2_io_validout64_15),
    .io_validout64_16(ingress2_io_validout64_16),
    .io_validout64_17(ingress2_io_validout64_17),
    .io_validout64_18(ingress2_io_validout64_18),
    .io_validout64_19(ingress2_io_validout64_19),
    .io_validout64_20(ingress2_io_validout64_20),
    .io_validout64_21(ingress2_io_validout64_21),
    .io_validout64_22(ingress2_io_validout64_22),
    .io_validout64_23(ingress2_io_validout64_23),
    .io_validout64_24(ingress2_io_validout64_24),
    .io_validout64_25(ingress2_io_validout64_25),
    .io_validout64_26(ingress2_io_validout64_26),
    .io_validout64_27(ingress2_io_validout64_27),
    .io_validout64_28(ingress2_io_validout64_28),
    .io_validout64_29(ingress2_io_validout64_29),
    .io_validout64_30(ingress2_io_validout64_30),
    .io_validout64_31(ingress2_io_validout64_31),
    .io_validout64_32(ingress2_io_validout64_32),
    .io_validout64_33(ingress2_io_validout64_33),
    .io_validout64_34(ingress2_io_validout64_34),
    .io_validout64_35(ingress2_io_validout64_35),
    .io_validout64_36(ingress2_io_validout64_36),
    .io_validout64_37(ingress2_io_validout64_37),
    .io_validout64_38(ingress2_io_validout64_38),
    .io_validout64_39(ingress2_io_validout64_39),
    .io_validout64_40(ingress2_io_validout64_40),
    .io_validout64_41(ingress2_io_validout64_41),
    .io_validout64_42(ingress2_io_validout64_42),
    .io_validout64_43(ingress2_io_validout64_43),
    .io_validout64_44(ingress2_io_validout64_44),
    .io_validout64_45(ingress2_io_validout64_45),
    .io_validout64_46(ingress2_io_validout64_46),
    .io_validout64_47(ingress2_io_validout64_47),
    .io_validout64_48(ingress2_io_validout64_48),
    .io_validout64_49(ingress2_io_validout64_49),
    .io_validout64_50(ingress2_io_validout64_50),
    .io_validout64_51(ingress2_io_validout64_51),
    .io_validout64_52(ingress2_io_validout64_52),
    .io_validout64_53(ingress2_io_validout64_53),
    .io_validout64_54(ingress2_io_validout64_54),
    .io_validout64_55(ingress2_io_validout64_55),
    .io_validout64_56(ingress2_io_validout64_56),
    .io_validout64_57(ingress2_io_validout64_57),
    .io_validout64_58(ingress2_io_validout64_58),
    .io_validout64_59(ingress2_io_validout64_59),
    .io_validout64_60(ingress2_io_validout64_60),
    .io_validout64_61(ingress2_io_validout64_61),
    .io_validout64_62(ingress2_io_validout64_62),
    .io_validout64_63(ingress2_io_validout64_63),
    .io_addrout(ingress2_io_addrout),
    .io_ctrl(ingress2_io_ctrl)
  );
  CLOSingress2 middle ( // @[BuildingBlockNew.scala 86:22]
    .clock(middle_clock),
    .io_in64_0(middle_io_in64_0),
    .io_in64_1(middle_io_in64_1),
    .io_in64_2(middle_io_in64_2),
    .io_in64_3(middle_io_in64_3),
    .io_in64_4(middle_io_in64_4),
    .io_in64_5(middle_io_in64_5),
    .io_in64_6(middle_io_in64_6),
    .io_in64_7(middle_io_in64_7),
    .io_in64_8(middle_io_in64_8),
    .io_in64_9(middle_io_in64_9),
    .io_in64_10(middle_io_in64_10),
    .io_in64_11(middle_io_in64_11),
    .io_in64_12(middle_io_in64_12),
    .io_in64_13(middle_io_in64_13),
    .io_in64_14(middle_io_in64_14),
    .io_in64_15(middle_io_in64_15),
    .io_in64_16(middle_io_in64_16),
    .io_in64_17(middle_io_in64_17),
    .io_in64_18(middle_io_in64_18),
    .io_in64_19(middle_io_in64_19),
    .io_in64_20(middle_io_in64_20),
    .io_in64_21(middle_io_in64_21),
    .io_in64_22(middle_io_in64_22),
    .io_in64_23(middle_io_in64_23),
    .io_in64_24(middle_io_in64_24),
    .io_in64_25(middle_io_in64_25),
    .io_in64_26(middle_io_in64_26),
    .io_in64_27(middle_io_in64_27),
    .io_in64_28(middle_io_in64_28),
    .io_in64_29(middle_io_in64_29),
    .io_in64_30(middle_io_in64_30),
    .io_in64_31(middle_io_in64_31),
    .io_in64_32(middle_io_in64_32),
    .io_in64_33(middle_io_in64_33),
    .io_in64_34(middle_io_in64_34),
    .io_in64_35(middle_io_in64_35),
    .io_in64_36(middle_io_in64_36),
    .io_in64_37(middle_io_in64_37),
    .io_in64_38(middle_io_in64_38),
    .io_in64_39(middle_io_in64_39),
    .io_in64_40(middle_io_in64_40),
    .io_in64_41(middle_io_in64_41),
    .io_in64_42(middle_io_in64_42),
    .io_in64_43(middle_io_in64_43),
    .io_in64_44(middle_io_in64_44),
    .io_in64_45(middle_io_in64_45),
    .io_in64_46(middle_io_in64_46),
    .io_in64_47(middle_io_in64_47),
    .io_in64_48(middle_io_in64_48),
    .io_in64_49(middle_io_in64_49),
    .io_in64_50(middle_io_in64_50),
    .io_in64_51(middle_io_in64_51),
    .io_in64_52(middle_io_in64_52),
    .io_in64_53(middle_io_in64_53),
    .io_in64_54(middle_io_in64_54),
    .io_in64_55(middle_io_in64_55),
    .io_in64_56(middle_io_in64_56),
    .io_in64_57(middle_io_in64_57),
    .io_in64_58(middle_io_in64_58),
    .io_in64_59(middle_io_in64_59),
    .io_in64_60(middle_io_in64_60),
    .io_in64_61(middle_io_in64_61),
    .io_in64_62(middle_io_in64_62),
    .io_in64_63(middle_io_in64_63),
    .io_validin64_0(middle_io_validin64_0),
    .io_validin64_1(middle_io_validin64_1),
    .io_validin64_2(middle_io_validin64_2),
    .io_validin64_3(middle_io_validin64_3),
    .io_validin64_4(middle_io_validin64_4),
    .io_validin64_5(middle_io_validin64_5),
    .io_validin64_6(middle_io_validin64_6),
    .io_validin64_7(middle_io_validin64_7),
    .io_validin64_8(middle_io_validin64_8),
    .io_validin64_9(middle_io_validin64_9),
    .io_validin64_10(middle_io_validin64_10),
    .io_validin64_11(middle_io_validin64_11),
    .io_validin64_12(middle_io_validin64_12),
    .io_validin64_13(middle_io_validin64_13),
    .io_validin64_14(middle_io_validin64_14),
    .io_validin64_15(middle_io_validin64_15),
    .io_validin64_16(middle_io_validin64_16),
    .io_validin64_17(middle_io_validin64_17),
    .io_validin64_18(middle_io_validin64_18),
    .io_validin64_19(middle_io_validin64_19),
    .io_validin64_20(middle_io_validin64_20),
    .io_validin64_21(middle_io_validin64_21),
    .io_validin64_22(middle_io_validin64_22),
    .io_validin64_23(middle_io_validin64_23),
    .io_validin64_24(middle_io_validin64_24),
    .io_validin64_25(middle_io_validin64_25),
    .io_validin64_26(middle_io_validin64_26),
    .io_validin64_27(middle_io_validin64_27),
    .io_validin64_28(middle_io_validin64_28),
    .io_validin64_29(middle_io_validin64_29),
    .io_validin64_30(middle_io_validin64_30),
    .io_validin64_31(middle_io_validin64_31),
    .io_validin64_32(middle_io_validin64_32),
    .io_validin64_33(middle_io_validin64_33),
    .io_validin64_34(middle_io_validin64_34),
    .io_validin64_35(middle_io_validin64_35),
    .io_validin64_36(middle_io_validin64_36),
    .io_validin64_37(middle_io_validin64_37),
    .io_validin64_38(middle_io_validin64_38),
    .io_validin64_39(middle_io_validin64_39),
    .io_validin64_40(middle_io_validin64_40),
    .io_validin64_41(middle_io_validin64_41),
    .io_validin64_42(middle_io_validin64_42),
    .io_validin64_43(middle_io_validin64_43),
    .io_validin64_44(middle_io_validin64_44),
    .io_validin64_45(middle_io_validin64_45),
    .io_validin64_46(middle_io_validin64_46),
    .io_validin64_47(middle_io_validin64_47),
    .io_validin64_48(middle_io_validin64_48),
    .io_validin64_49(middle_io_validin64_49),
    .io_validin64_50(middle_io_validin64_50),
    .io_validin64_51(middle_io_validin64_51),
    .io_validin64_52(middle_io_validin64_52),
    .io_validin64_53(middle_io_validin64_53),
    .io_validin64_54(middle_io_validin64_54),
    .io_validin64_55(middle_io_validin64_55),
    .io_validin64_56(middle_io_validin64_56),
    .io_validin64_57(middle_io_validin64_57),
    .io_validin64_58(middle_io_validin64_58),
    .io_validin64_59(middle_io_validin64_59),
    .io_validin64_60(middle_io_validin64_60),
    .io_validin64_61(middle_io_validin64_61),
    .io_validin64_62(middle_io_validin64_62),
    .io_validin64_63(middle_io_validin64_63),
    .io_addrin(middle_io_addrin),
    .io_out64_0(middle_io_out64_0),
    .io_out64_1(middle_io_out64_1),
    .io_out64_2(middle_io_out64_2),
    .io_out64_3(middle_io_out64_3),
    .io_out64_4(middle_io_out64_4),
    .io_out64_5(middle_io_out64_5),
    .io_out64_6(middle_io_out64_6),
    .io_out64_7(middle_io_out64_7),
    .io_out64_8(middle_io_out64_8),
    .io_out64_9(middle_io_out64_9),
    .io_out64_10(middle_io_out64_10),
    .io_out64_11(middle_io_out64_11),
    .io_out64_12(middle_io_out64_12),
    .io_out64_13(middle_io_out64_13),
    .io_out64_14(middle_io_out64_14),
    .io_out64_15(middle_io_out64_15),
    .io_out64_16(middle_io_out64_16),
    .io_out64_17(middle_io_out64_17),
    .io_out64_18(middle_io_out64_18),
    .io_out64_19(middle_io_out64_19),
    .io_out64_20(middle_io_out64_20),
    .io_out64_21(middle_io_out64_21),
    .io_out64_22(middle_io_out64_22),
    .io_out64_23(middle_io_out64_23),
    .io_out64_24(middle_io_out64_24),
    .io_out64_25(middle_io_out64_25),
    .io_out64_26(middle_io_out64_26),
    .io_out64_27(middle_io_out64_27),
    .io_out64_28(middle_io_out64_28),
    .io_out64_29(middle_io_out64_29),
    .io_out64_30(middle_io_out64_30),
    .io_out64_31(middle_io_out64_31),
    .io_out64_32(middle_io_out64_32),
    .io_out64_33(middle_io_out64_33),
    .io_out64_34(middle_io_out64_34),
    .io_out64_35(middle_io_out64_35),
    .io_out64_36(middle_io_out64_36),
    .io_out64_37(middle_io_out64_37),
    .io_out64_38(middle_io_out64_38),
    .io_out64_39(middle_io_out64_39),
    .io_out64_40(middle_io_out64_40),
    .io_out64_41(middle_io_out64_41),
    .io_out64_42(middle_io_out64_42),
    .io_out64_43(middle_io_out64_43),
    .io_out64_44(middle_io_out64_44),
    .io_out64_45(middle_io_out64_45),
    .io_out64_46(middle_io_out64_46),
    .io_out64_47(middle_io_out64_47),
    .io_out64_48(middle_io_out64_48),
    .io_out64_49(middle_io_out64_49),
    .io_out64_50(middle_io_out64_50),
    .io_out64_51(middle_io_out64_51),
    .io_out64_52(middle_io_out64_52),
    .io_out64_53(middle_io_out64_53),
    .io_out64_54(middle_io_out64_54),
    .io_out64_55(middle_io_out64_55),
    .io_out64_56(middle_io_out64_56),
    .io_out64_57(middle_io_out64_57),
    .io_out64_58(middle_io_out64_58),
    .io_out64_59(middle_io_out64_59),
    .io_out64_60(middle_io_out64_60),
    .io_out64_61(middle_io_out64_61),
    .io_out64_62(middle_io_out64_62),
    .io_out64_63(middle_io_out64_63),
    .io_validout64_0(middle_io_validout64_0),
    .io_validout64_1(middle_io_validout64_1),
    .io_validout64_2(middle_io_validout64_2),
    .io_validout64_3(middle_io_validout64_3),
    .io_validout64_4(middle_io_validout64_4),
    .io_validout64_5(middle_io_validout64_5),
    .io_validout64_6(middle_io_validout64_6),
    .io_validout64_7(middle_io_validout64_7),
    .io_validout64_8(middle_io_validout64_8),
    .io_validout64_9(middle_io_validout64_9),
    .io_validout64_10(middle_io_validout64_10),
    .io_validout64_11(middle_io_validout64_11),
    .io_validout64_12(middle_io_validout64_12),
    .io_validout64_13(middle_io_validout64_13),
    .io_validout64_14(middle_io_validout64_14),
    .io_validout64_15(middle_io_validout64_15),
    .io_validout64_16(middle_io_validout64_16),
    .io_validout64_17(middle_io_validout64_17),
    .io_validout64_18(middle_io_validout64_18),
    .io_validout64_19(middle_io_validout64_19),
    .io_validout64_20(middle_io_validout64_20),
    .io_validout64_21(middle_io_validout64_21),
    .io_validout64_22(middle_io_validout64_22),
    .io_validout64_23(middle_io_validout64_23),
    .io_validout64_24(middle_io_validout64_24),
    .io_validout64_25(middle_io_validout64_25),
    .io_validout64_26(middle_io_validout64_26),
    .io_validout64_27(middle_io_validout64_27),
    .io_validout64_28(middle_io_validout64_28),
    .io_validout64_29(middle_io_validout64_29),
    .io_validout64_30(middle_io_validout64_30),
    .io_validout64_31(middle_io_validout64_31),
    .io_validout64_32(middle_io_validout64_32),
    .io_validout64_33(middle_io_validout64_33),
    .io_validout64_34(middle_io_validout64_34),
    .io_validout64_35(middle_io_validout64_35),
    .io_validout64_36(middle_io_validout64_36),
    .io_validout64_37(middle_io_validout64_37),
    .io_validout64_38(middle_io_validout64_38),
    .io_validout64_39(middle_io_validout64_39),
    .io_validout64_40(middle_io_validout64_40),
    .io_validout64_41(middle_io_validout64_41),
    .io_validout64_42(middle_io_validout64_42),
    .io_validout64_43(middle_io_validout64_43),
    .io_validout64_44(middle_io_validout64_44),
    .io_validout64_45(middle_io_validout64_45),
    .io_validout64_46(middle_io_validout64_46),
    .io_validout64_47(middle_io_validout64_47),
    .io_validout64_48(middle_io_validout64_48),
    .io_validout64_49(middle_io_validout64_49),
    .io_validout64_50(middle_io_validout64_50),
    .io_validout64_51(middle_io_validout64_51),
    .io_validout64_52(middle_io_validout64_52),
    .io_validout64_53(middle_io_validout64_53),
    .io_validout64_54(middle_io_validout64_54),
    .io_validout64_55(middle_io_validout64_55),
    .io_validout64_56(middle_io_validout64_56),
    .io_validout64_57(middle_io_validout64_57),
    .io_validout64_58(middle_io_validout64_58),
    .io_validout64_59(middle_io_validout64_59),
    .io_validout64_60(middle_io_validout64_60),
    .io_validout64_61(middle_io_validout64_61),
    .io_validout64_62(middle_io_validout64_62),
    .io_validout64_63(middle_io_validout64_63),
    .io_addrout(middle_io_addrout),
    .io_ctrl(middle_io_ctrl)
  );
  CLOSegress1 egress1 ( // @[BuildingBlockNew.scala 87:23]
    .clock(egress1_clock),
    .io_in64_0(egress1_io_in64_0),
    .io_in64_1(egress1_io_in64_1),
    .io_in64_2(egress1_io_in64_2),
    .io_in64_3(egress1_io_in64_3),
    .io_in64_4(egress1_io_in64_4),
    .io_in64_5(egress1_io_in64_5),
    .io_in64_6(egress1_io_in64_6),
    .io_in64_7(egress1_io_in64_7),
    .io_in64_8(egress1_io_in64_8),
    .io_in64_9(egress1_io_in64_9),
    .io_in64_10(egress1_io_in64_10),
    .io_in64_11(egress1_io_in64_11),
    .io_in64_12(egress1_io_in64_12),
    .io_in64_13(egress1_io_in64_13),
    .io_in64_14(egress1_io_in64_14),
    .io_in64_15(egress1_io_in64_15),
    .io_in64_16(egress1_io_in64_16),
    .io_in64_17(egress1_io_in64_17),
    .io_in64_18(egress1_io_in64_18),
    .io_in64_19(egress1_io_in64_19),
    .io_in64_20(egress1_io_in64_20),
    .io_in64_21(egress1_io_in64_21),
    .io_in64_22(egress1_io_in64_22),
    .io_in64_23(egress1_io_in64_23),
    .io_in64_24(egress1_io_in64_24),
    .io_in64_25(egress1_io_in64_25),
    .io_in64_26(egress1_io_in64_26),
    .io_in64_27(egress1_io_in64_27),
    .io_in64_28(egress1_io_in64_28),
    .io_in64_29(egress1_io_in64_29),
    .io_in64_30(egress1_io_in64_30),
    .io_in64_31(egress1_io_in64_31),
    .io_in64_32(egress1_io_in64_32),
    .io_in64_33(egress1_io_in64_33),
    .io_in64_34(egress1_io_in64_34),
    .io_in64_35(egress1_io_in64_35),
    .io_in64_36(egress1_io_in64_36),
    .io_in64_37(egress1_io_in64_37),
    .io_in64_38(egress1_io_in64_38),
    .io_in64_39(egress1_io_in64_39),
    .io_in64_40(egress1_io_in64_40),
    .io_in64_41(egress1_io_in64_41),
    .io_in64_42(egress1_io_in64_42),
    .io_in64_43(egress1_io_in64_43),
    .io_in64_44(egress1_io_in64_44),
    .io_in64_45(egress1_io_in64_45),
    .io_in64_46(egress1_io_in64_46),
    .io_in64_47(egress1_io_in64_47),
    .io_in64_48(egress1_io_in64_48),
    .io_in64_49(egress1_io_in64_49),
    .io_in64_50(egress1_io_in64_50),
    .io_in64_51(egress1_io_in64_51),
    .io_in64_52(egress1_io_in64_52),
    .io_in64_53(egress1_io_in64_53),
    .io_in64_54(egress1_io_in64_54),
    .io_in64_55(egress1_io_in64_55),
    .io_in64_56(egress1_io_in64_56),
    .io_in64_57(egress1_io_in64_57),
    .io_in64_58(egress1_io_in64_58),
    .io_in64_59(egress1_io_in64_59),
    .io_in64_60(egress1_io_in64_60),
    .io_in64_61(egress1_io_in64_61),
    .io_in64_62(egress1_io_in64_62),
    .io_in64_63(egress1_io_in64_63),
    .io_validin64_0(egress1_io_validin64_0),
    .io_validin64_1(egress1_io_validin64_1),
    .io_validin64_2(egress1_io_validin64_2),
    .io_validin64_3(egress1_io_validin64_3),
    .io_validin64_4(egress1_io_validin64_4),
    .io_validin64_5(egress1_io_validin64_5),
    .io_validin64_6(egress1_io_validin64_6),
    .io_validin64_7(egress1_io_validin64_7),
    .io_validin64_8(egress1_io_validin64_8),
    .io_validin64_9(egress1_io_validin64_9),
    .io_validin64_10(egress1_io_validin64_10),
    .io_validin64_11(egress1_io_validin64_11),
    .io_validin64_12(egress1_io_validin64_12),
    .io_validin64_13(egress1_io_validin64_13),
    .io_validin64_14(egress1_io_validin64_14),
    .io_validin64_15(egress1_io_validin64_15),
    .io_validin64_16(egress1_io_validin64_16),
    .io_validin64_17(egress1_io_validin64_17),
    .io_validin64_18(egress1_io_validin64_18),
    .io_validin64_19(egress1_io_validin64_19),
    .io_validin64_20(egress1_io_validin64_20),
    .io_validin64_21(egress1_io_validin64_21),
    .io_validin64_22(egress1_io_validin64_22),
    .io_validin64_23(egress1_io_validin64_23),
    .io_validin64_24(egress1_io_validin64_24),
    .io_validin64_25(egress1_io_validin64_25),
    .io_validin64_26(egress1_io_validin64_26),
    .io_validin64_27(egress1_io_validin64_27),
    .io_validin64_28(egress1_io_validin64_28),
    .io_validin64_29(egress1_io_validin64_29),
    .io_validin64_30(egress1_io_validin64_30),
    .io_validin64_31(egress1_io_validin64_31),
    .io_validin64_32(egress1_io_validin64_32),
    .io_validin64_33(egress1_io_validin64_33),
    .io_validin64_34(egress1_io_validin64_34),
    .io_validin64_35(egress1_io_validin64_35),
    .io_validin64_36(egress1_io_validin64_36),
    .io_validin64_37(egress1_io_validin64_37),
    .io_validin64_38(egress1_io_validin64_38),
    .io_validin64_39(egress1_io_validin64_39),
    .io_validin64_40(egress1_io_validin64_40),
    .io_validin64_41(egress1_io_validin64_41),
    .io_validin64_42(egress1_io_validin64_42),
    .io_validin64_43(egress1_io_validin64_43),
    .io_validin64_44(egress1_io_validin64_44),
    .io_validin64_45(egress1_io_validin64_45),
    .io_validin64_46(egress1_io_validin64_46),
    .io_validin64_47(egress1_io_validin64_47),
    .io_validin64_48(egress1_io_validin64_48),
    .io_validin64_49(egress1_io_validin64_49),
    .io_validin64_50(egress1_io_validin64_50),
    .io_validin64_51(egress1_io_validin64_51),
    .io_validin64_52(egress1_io_validin64_52),
    .io_validin64_53(egress1_io_validin64_53),
    .io_validin64_54(egress1_io_validin64_54),
    .io_validin64_55(egress1_io_validin64_55),
    .io_validin64_56(egress1_io_validin64_56),
    .io_validin64_57(egress1_io_validin64_57),
    .io_validin64_58(egress1_io_validin64_58),
    .io_validin64_59(egress1_io_validin64_59),
    .io_validin64_60(egress1_io_validin64_60),
    .io_validin64_61(egress1_io_validin64_61),
    .io_validin64_62(egress1_io_validin64_62),
    .io_validin64_63(egress1_io_validin64_63),
    .io_addrin(egress1_io_addrin),
    .io_out64_0(egress1_io_out64_0),
    .io_out64_1(egress1_io_out64_1),
    .io_out64_2(egress1_io_out64_2),
    .io_out64_3(egress1_io_out64_3),
    .io_out64_4(egress1_io_out64_4),
    .io_out64_5(egress1_io_out64_5),
    .io_out64_6(egress1_io_out64_6),
    .io_out64_7(egress1_io_out64_7),
    .io_out64_8(egress1_io_out64_8),
    .io_out64_9(egress1_io_out64_9),
    .io_out64_10(egress1_io_out64_10),
    .io_out64_11(egress1_io_out64_11),
    .io_out64_12(egress1_io_out64_12),
    .io_out64_13(egress1_io_out64_13),
    .io_out64_14(egress1_io_out64_14),
    .io_out64_15(egress1_io_out64_15),
    .io_out64_16(egress1_io_out64_16),
    .io_out64_17(egress1_io_out64_17),
    .io_out64_18(egress1_io_out64_18),
    .io_out64_19(egress1_io_out64_19),
    .io_out64_20(egress1_io_out64_20),
    .io_out64_21(egress1_io_out64_21),
    .io_out64_22(egress1_io_out64_22),
    .io_out64_23(egress1_io_out64_23),
    .io_out64_24(egress1_io_out64_24),
    .io_out64_25(egress1_io_out64_25),
    .io_out64_26(egress1_io_out64_26),
    .io_out64_27(egress1_io_out64_27),
    .io_out64_28(egress1_io_out64_28),
    .io_out64_29(egress1_io_out64_29),
    .io_out64_30(egress1_io_out64_30),
    .io_out64_31(egress1_io_out64_31),
    .io_out64_32(egress1_io_out64_32),
    .io_out64_33(egress1_io_out64_33),
    .io_out64_34(egress1_io_out64_34),
    .io_out64_35(egress1_io_out64_35),
    .io_out64_36(egress1_io_out64_36),
    .io_out64_37(egress1_io_out64_37),
    .io_out64_38(egress1_io_out64_38),
    .io_out64_39(egress1_io_out64_39),
    .io_out64_40(egress1_io_out64_40),
    .io_out64_41(egress1_io_out64_41),
    .io_out64_42(egress1_io_out64_42),
    .io_out64_43(egress1_io_out64_43),
    .io_out64_44(egress1_io_out64_44),
    .io_out64_45(egress1_io_out64_45),
    .io_out64_46(egress1_io_out64_46),
    .io_out64_47(egress1_io_out64_47),
    .io_out64_48(egress1_io_out64_48),
    .io_out64_49(egress1_io_out64_49),
    .io_out64_50(egress1_io_out64_50),
    .io_out64_51(egress1_io_out64_51),
    .io_out64_52(egress1_io_out64_52),
    .io_out64_53(egress1_io_out64_53),
    .io_out64_54(egress1_io_out64_54),
    .io_out64_55(egress1_io_out64_55),
    .io_out64_56(egress1_io_out64_56),
    .io_out64_57(egress1_io_out64_57),
    .io_out64_58(egress1_io_out64_58),
    .io_out64_59(egress1_io_out64_59),
    .io_out64_60(egress1_io_out64_60),
    .io_out64_61(egress1_io_out64_61),
    .io_out64_62(egress1_io_out64_62),
    .io_out64_63(egress1_io_out64_63),
    .io_validout64_0(egress1_io_validout64_0),
    .io_validout64_1(egress1_io_validout64_1),
    .io_validout64_2(egress1_io_validout64_2),
    .io_validout64_3(egress1_io_validout64_3),
    .io_validout64_4(egress1_io_validout64_4),
    .io_validout64_5(egress1_io_validout64_5),
    .io_validout64_6(egress1_io_validout64_6),
    .io_validout64_7(egress1_io_validout64_7),
    .io_validout64_8(egress1_io_validout64_8),
    .io_validout64_9(egress1_io_validout64_9),
    .io_validout64_10(egress1_io_validout64_10),
    .io_validout64_11(egress1_io_validout64_11),
    .io_validout64_12(egress1_io_validout64_12),
    .io_validout64_13(egress1_io_validout64_13),
    .io_validout64_14(egress1_io_validout64_14),
    .io_validout64_15(egress1_io_validout64_15),
    .io_validout64_16(egress1_io_validout64_16),
    .io_validout64_17(egress1_io_validout64_17),
    .io_validout64_18(egress1_io_validout64_18),
    .io_validout64_19(egress1_io_validout64_19),
    .io_validout64_20(egress1_io_validout64_20),
    .io_validout64_21(egress1_io_validout64_21),
    .io_validout64_22(egress1_io_validout64_22),
    .io_validout64_23(egress1_io_validout64_23),
    .io_validout64_24(egress1_io_validout64_24),
    .io_validout64_25(egress1_io_validout64_25),
    .io_validout64_26(egress1_io_validout64_26),
    .io_validout64_27(egress1_io_validout64_27),
    .io_validout64_28(egress1_io_validout64_28),
    .io_validout64_29(egress1_io_validout64_29),
    .io_validout64_30(egress1_io_validout64_30),
    .io_validout64_31(egress1_io_validout64_31),
    .io_validout64_32(egress1_io_validout64_32),
    .io_validout64_33(egress1_io_validout64_33),
    .io_validout64_34(egress1_io_validout64_34),
    .io_validout64_35(egress1_io_validout64_35),
    .io_validout64_36(egress1_io_validout64_36),
    .io_validout64_37(egress1_io_validout64_37),
    .io_validout64_38(egress1_io_validout64_38),
    .io_validout64_39(egress1_io_validout64_39),
    .io_validout64_40(egress1_io_validout64_40),
    .io_validout64_41(egress1_io_validout64_41),
    .io_validout64_42(egress1_io_validout64_42),
    .io_validout64_43(egress1_io_validout64_43),
    .io_validout64_44(egress1_io_validout64_44),
    .io_validout64_45(egress1_io_validout64_45),
    .io_validout64_46(egress1_io_validout64_46),
    .io_validout64_47(egress1_io_validout64_47),
    .io_validout64_48(egress1_io_validout64_48),
    .io_validout64_49(egress1_io_validout64_49),
    .io_validout64_50(egress1_io_validout64_50),
    .io_validout64_51(egress1_io_validout64_51),
    .io_validout64_52(egress1_io_validout64_52),
    .io_validout64_53(egress1_io_validout64_53),
    .io_validout64_54(egress1_io_validout64_54),
    .io_validout64_55(egress1_io_validout64_55),
    .io_validout64_56(egress1_io_validout64_56),
    .io_validout64_57(egress1_io_validout64_57),
    .io_validout64_58(egress1_io_validout64_58),
    .io_validout64_59(egress1_io_validout64_59),
    .io_validout64_60(egress1_io_validout64_60),
    .io_validout64_61(egress1_io_validout64_61),
    .io_validout64_62(egress1_io_validout64_62),
    .io_validout64_63(egress1_io_validout64_63),
    .io_addrout(egress1_io_addrout),
    .io_ctrl(egress1_io_ctrl)
  );
  CLOSegress2 egress2 ( // @[BuildingBlockNew.scala 88:23]
    .clock(egress2_clock),
    .io_in64_0(egress2_io_in64_0),
    .io_in64_1(egress2_io_in64_1),
    .io_in64_2(egress2_io_in64_2),
    .io_in64_3(egress2_io_in64_3),
    .io_in64_4(egress2_io_in64_4),
    .io_in64_5(egress2_io_in64_5),
    .io_in64_6(egress2_io_in64_6),
    .io_in64_7(egress2_io_in64_7),
    .io_in64_8(egress2_io_in64_8),
    .io_in64_9(egress2_io_in64_9),
    .io_in64_10(egress2_io_in64_10),
    .io_in64_11(egress2_io_in64_11),
    .io_in64_12(egress2_io_in64_12),
    .io_in64_13(egress2_io_in64_13),
    .io_in64_14(egress2_io_in64_14),
    .io_in64_15(egress2_io_in64_15),
    .io_in64_16(egress2_io_in64_16),
    .io_in64_17(egress2_io_in64_17),
    .io_in64_18(egress2_io_in64_18),
    .io_in64_19(egress2_io_in64_19),
    .io_in64_20(egress2_io_in64_20),
    .io_in64_21(egress2_io_in64_21),
    .io_in64_22(egress2_io_in64_22),
    .io_in64_23(egress2_io_in64_23),
    .io_in64_24(egress2_io_in64_24),
    .io_in64_25(egress2_io_in64_25),
    .io_in64_26(egress2_io_in64_26),
    .io_in64_27(egress2_io_in64_27),
    .io_in64_28(egress2_io_in64_28),
    .io_in64_29(egress2_io_in64_29),
    .io_in64_30(egress2_io_in64_30),
    .io_in64_31(egress2_io_in64_31),
    .io_in64_32(egress2_io_in64_32),
    .io_in64_33(egress2_io_in64_33),
    .io_in64_34(egress2_io_in64_34),
    .io_in64_35(egress2_io_in64_35),
    .io_in64_36(egress2_io_in64_36),
    .io_in64_37(egress2_io_in64_37),
    .io_in64_38(egress2_io_in64_38),
    .io_in64_39(egress2_io_in64_39),
    .io_in64_40(egress2_io_in64_40),
    .io_in64_41(egress2_io_in64_41),
    .io_in64_42(egress2_io_in64_42),
    .io_in64_43(egress2_io_in64_43),
    .io_in64_44(egress2_io_in64_44),
    .io_in64_45(egress2_io_in64_45),
    .io_in64_46(egress2_io_in64_46),
    .io_in64_47(egress2_io_in64_47),
    .io_in64_48(egress2_io_in64_48),
    .io_in64_49(egress2_io_in64_49),
    .io_in64_50(egress2_io_in64_50),
    .io_in64_51(egress2_io_in64_51),
    .io_in64_52(egress2_io_in64_52),
    .io_in64_53(egress2_io_in64_53),
    .io_in64_54(egress2_io_in64_54),
    .io_in64_55(egress2_io_in64_55),
    .io_in64_56(egress2_io_in64_56),
    .io_in64_57(egress2_io_in64_57),
    .io_in64_58(egress2_io_in64_58),
    .io_in64_59(egress2_io_in64_59),
    .io_in64_60(egress2_io_in64_60),
    .io_in64_61(egress2_io_in64_61),
    .io_in64_62(egress2_io_in64_62),
    .io_in64_63(egress2_io_in64_63),
    .io_validin64_0(egress2_io_validin64_0),
    .io_validin64_1(egress2_io_validin64_1),
    .io_validin64_2(egress2_io_validin64_2),
    .io_validin64_3(egress2_io_validin64_3),
    .io_validin64_4(egress2_io_validin64_4),
    .io_validin64_5(egress2_io_validin64_5),
    .io_validin64_6(egress2_io_validin64_6),
    .io_validin64_7(egress2_io_validin64_7),
    .io_validin64_8(egress2_io_validin64_8),
    .io_validin64_9(egress2_io_validin64_9),
    .io_validin64_10(egress2_io_validin64_10),
    .io_validin64_11(egress2_io_validin64_11),
    .io_validin64_12(egress2_io_validin64_12),
    .io_validin64_13(egress2_io_validin64_13),
    .io_validin64_14(egress2_io_validin64_14),
    .io_validin64_15(egress2_io_validin64_15),
    .io_validin64_16(egress2_io_validin64_16),
    .io_validin64_17(egress2_io_validin64_17),
    .io_validin64_18(egress2_io_validin64_18),
    .io_validin64_19(egress2_io_validin64_19),
    .io_validin64_20(egress2_io_validin64_20),
    .io_validin64_21(egress2_io_validin64_21),
    .io_validin64_22(egress2_io_validin64_22),
    .io_validin64_23(egress2_io_validin64_23),
    .io_validin64_24(egress2_io_validin64_24),
    .io_validin64_25(egress2_io_validin64_25),
    .io_validin64_26(egress2_io_validin64_26),
    .io_validin64_27(egress2_io_validin64_27),
    .io_validin64_28(egress2_io_validin64_28),
    .io_validin64_29(egress2_io_validin64_29),
    .io_validin64_30(egress2_io_validin64_30),
    .io_validin64_31(egress2_io_validin64_31),
    .io_validin64_32(egress2_io_validin64_32),
    .io_validin64_33(egress2_io_validin64_33),
    .io_validin64_34(egress2_io_validin64_34),
    .io_validin64_35(egress2_io_validin64_35),
    .io_validin64_36(egress2_io_validin64_36),
    .io_validin64_37(egress2_io_validin64_37),
    .io_validin64_38(egress2_io_validin64_38),
    .io_validin64_39(egress2_io_validin64_39),
    .io_validin64_40(egress2_io_validin64_40),
    .io_validin64_41(egress2_io_validin64_41),
    .io_validin64_42(egress2_io_validin64_42),
    .io_validin64_43(egress2_io_validin64_43),
    .io_validin64_44(egress2_io_validin64_44),
    .io_validin64_45(egress2_io_validin64_45),
    .io_validin64_46(egress2_io_validin64_46),
    .io_validin64_47(egress2_io_validin64_47),
    .io_validin64_48(egress2_io_validin64_48),
    .io_validin64_49(egress2_io_validin64_49),
    .io_validin64_50(egress2_io_validin64_50),
    .io_validin64_51(egress2_io_validin64_51),
    .io_validin64_52(egress2_io_validin64_52),
    .io_validin64_53(egress2_io_validin64_53),
    .io_validin64_54(egress2_io_validin64_54),
    .io_validin64_55(egress2_io_validin64_55),
    .io_validin64_56(egress2_io_validin64_56),
    .io_validin64_57(egress2_io_validin64_57),
    .io_validin64_58(egress2_io_validin64_58),
    .io_validin64_59(egress2_io_validin64_59),
    .io_validin64_60(egress2_io_validin64_60),
    .io_validin64_61(egress2_io_validin64_61),
    .io_validin64_62(egress2_io_validin64_62),
    .io_validin64_63(egress2_io_validin64_63),
    .io_addrin(egress2_io_addrin),
    .io_out64_0(egress2_io_out64_0),
    .io_out64_1(egress2_io_out64_1),
    .io_out64_2(egress2_io_out64_2),
    .io_out64_3(egress2_io_out64_3),
    .io_out64_4(egress2_io_out64_4),
    .io_out64_5(egress2_io_out64_5),
    .io_out64_6(egress2_io_out64_6),
    .io_out64_7(egress2_io_out64_7),
    .io_out64_8(egress2_io_out64_8),
    .io_out64_9(egress2_io_out64_9),
    .io_out64_10(egress2_io_out64_10),
    .io_out64_11(egress2_io_out64_11),
    .io_out64_12(egress2_io_out64_12),
    .io_out64_13(egress2_io_out64_13),
    .io_out64_14(egress2_io_out64_14),
    .io_out64_15(egress2_io_out64_15),
    .io_out64_16(egress2_io_out64_16),
    .io_out64_17(egress2_io_out64_17),
    .io_out64_18(egress2_io_out64_18),
    .io_out64_19(egress2_io_out64_19),
    .io_out64_20(egress2_io_out64_20),
    .io_out64_21(egress2_io_out64_21),
    .io_out64_22(egress2_io_out64_22),
    .io_out64_23(egress2_io_out64_23),
    .io_out64_24(egress2_io_out64_24),
    .io_out64_25(egress2_io_out64_25),
    .io_out64_26(egress2_io_out64_26),
    .io_out64_27(egress2_io_out64_27),
    .io_out64_28(egress2_io_out64_28),
    .io_out64_29(egress2_io_out64_29),
    .io_out64_30(egress2_io_out64_30),
    .io_out64_31(egress2_io_out64_31),
    .io_out64_32(egress2_io_out64_32),
    .io_out64_33(egress2_io_out64_33),
    .io_out64_34(egress2_io_out64_34),
    .io_out64_35(egress2_io_out64_35),
    .io_out64_36(egress2_io_out64_36),
    .io_out64_37(egress2_io_out64_37),
    .io_out64_38(egress2_io_out64_38),
    .io_out64_39(egress2_io_out64_39),
    .io_out64_40(egress2_io_out64_40),
    .io_out64_41(egress2_io_out64_41),
    .io_out64_42(egress2_io_out64_42),
    .io_out64_43(egress2_io_out64_43),
    .io_out64_44(egress2_io_out64_44),
    .io_out64_45(egress2_io_out64_45),
    .io_out64_46(egress2_io_out64_46),
    .io_out64_47(egress2_io_out64_47),
    .io_out64_48(egress2_io_out64_48),
    .io_out64_49(egress2_io_out64_49),
    .io_out64_50(egress2_io_out64_50),
    .io_out64_51(egress2_io_out64_51),
    .io_out64_52(egress2_io_out64_52),
    .io_out64_53(egress2_io_out64_53),
    .io_out64_54(egress2_io_out64_54),
    .io_out64_55(egress2_io_out64_55),
    .io_out64_56(egress2_io_out64_56),
    .io_out64_57(egress2_io_out64_57),
    .io_out64_58(egress2_io_out64_58),
    .io_out64_59(egress2_io_out64_59),
    .io_out64_60(egress2_io_out64_60),
    .io_out64_61(egress2_io_out64_61),
    .io_out64_62(egress2_io_out64_62),
    .io_out64_63(egress2_io_out64_63),
    .io_validout64_0(egress2_io_validout64_0),
    .io_validout64_1(egress2_io_validout64_1),
    .io_validout64_2(egress2_io_validout64_2),
    .io_validout64_3(egress2_io_validout64_3),
    .io_validout64_4(egress2_io_validout64_4),
    .io_validout64_5(egress2_io_validout64_5),
    .io_validout64_6(egress2_io_validout64_6),
    .io_validout64_7(egress2_io_validout64_7),
    .io_validout64_8(egress2_io_validout64_8),
    .io_validout64_9(egress2_io_validout64_9),
    .io_validout64_10(egress2_io_validout64_10),
    .io_validout64_11(egress2_io_validout64_11),
    .io_validout64_12(egress2_io_validout64_12),
    .io_validout64_13(egress2_io_validout64_13),
    .io_validout64_14(egress2_io_validout64_14),
    .io_validout64_15(egress2_io_validout64_15),
    .io_validout64_16(egress2_io_validout64_16),
    .io_validout64_17(egress2_io_validout64_17),
    .io_validout64_18(egress2_io_validout64_18),
    .io_validout64_19(egress2_io_validout64_19),
    .io_validout64_20(egress2_io_validout64_20),
    .io_validout64_21(egress2_io_validout64_21),
    .io_validout64_22(egress2_io_validout64_22),
    .io_validout64_23(egress2_io_validout64_23),
    .io_validout64_24(egress2_io_validout64_24),
    .io_validout64_25(egress2_io_validout64_25),
    .io_validout64_26(egress2_io_validout64_26),
    .io_validout64_27(egress2_io_validout64_27),
    .io_validout64_28(egress2_io_validout64_28),
    .io_validout64_29(egress2_io_validout64_29),
    .io_validout64_30(egress2_io_validout64_30),
    .io_validout64_31(egress2_io_validout64_31),
    .io_validout64_32(egress2_io_validout64_32),
    .io_validout64_33(egress2_io_validout64_33),
    .io_validout64_34(egress2_io_validout64_34),
    .io_validout64_35(egress2_io_validout64_35),
    .io_validout64_36(egress2_io_validout64_36),
    .io_validout64_37(egress2_io_validout64_37),
    .io_validout64_38(egress2_io_validout64_38),
    .io_validout64_39(egress2_io_validout64_39),
    .io_validout64_40(egress2_io_validout64_40),
    .io_validout64_41(egress2_io_validout64_41),
    .io_validout64_42(egress2_io_validout64_42),
    .io_validout64_43(egress2_io_validout64_43),
    .io_validout64_44(egress2_io_validout64_44),
    .io_validout64_45(egress2_io_validout64_45),
    .io_validout64_46(egress2_io_validout64_46),
    .io_validout64_47(egress2_io_validout64_47),
    .io_validout64_48(egress2_io_validout64_48),
    .io_validout64_49(egress2_io_validout64_49),
    .io_validout64_50(egress2_io_validout64_50),
    .io_validout64_51(egress2_io_validout64_51),
    .io_validout64_52(egress2_io_validout64_52),
    .io_validout64_53(egress2_io_validout64_53),
    .io_validout64_54(egress2_io_validout64_54),
    .io_validout64_55(egress2_io_validout64_55),
    .io_validout64_56(egress2_io_validout64_56),
    .io_validout64_57(egress2_io_validout64_57),
    .io_validout64_58(egress2_io_validout64_58),
    .io_validout64_59(egress2_io_validout64_59),
    .io_validout64_60(egress2_io_validout64_60),
    .io_validout64_61(egress2_io_validout64_61),
    .io_validout64_62(egress2_io_validout64_62),
    .io_validout64_63(egress2_io_validout64_63),
    .io_addrout(egress2_io_addrout),
    .io_ctrl(egress2_io_ctrl)
  );
  assign Mem1_instr1_MPORT_addr = Mem1_instr1_MPORT_addr_pipe_0;
  assign Mem1_instr1_MPORT_data = Mem1[Mem1_instr1_MPORT_addr]; // @[BuildingBlockNew.scala 33:25]
  assign Mem1_MPORT_data = io_wr_instr_mem1;
  assign Mem1_MPORT_addr = io_wr_en_mem1 ? wrAddr1 : PC1;
  assign Mem1_MPORT_mask = 1'h1;
  assign Mem1_MPORT_en = io_wr_en_mem1;
  assign Mem2_instr2_MPORT_addr = Mem2_instr2_MPORT_addr_pipe_0;
  assign Mem2_instr2_MPORT_data = Mem2[Mem2_instr2_MPORT_addr]; // @[BuildingBlockNew.scala 34:25]
  assign Mem2_MPORT_1_data = io_wr_instr_mem2;
  assign Mem2_MPORT_1_addr = io_wr_en_mem2 ? wrAddr2 : PC2;
  assign Mem2_MPORT_1_mask = 1'h1;
  assign Mem2_MPORT_1_en = io_wr_en_mem2;
  assign Mem3_instr3_MPORT_addr = Mem3_instr3_MPORT_addr_pipe_0;
  assign Mem3_instr3_MPORT_data = Mem3[Mem3_instr3_MPORT_addr]; // @[BuildingBlockNew.scala 35:25]
  assign Mem3_MPORT_2_data = io_wr_instr_mem3;
  assign Mem3_MPORT_2_addr = io_wr_en_mem3 ? wrAddr3 : PC3;
  assign Mem3_MPORT_2_mask = 1'h1;
  assign Mem3_MPORT_2_en = io_wr_en_mem3;
  assign Mem4_instr4_MPORT_addr = Mem4_instr4_MPORT_addr_pipe_0;
  assign Mem4_instr4_MPORT_data = Mem4[Mem4_instr4_MPORT_addr]; // @[BuildingBlockNew.scala 36:25]
  assign Mem4_MPORT_3_data = io_wr_instr_mem4;
  assign Mem4_MPORT_3_addr = io_wr_en_mem4 ? wrAddr4 : PC4;
  assign Mem4_MPORT_3_mask = 1'h1;
  assign Mem4_MPORT_3_en = io_wr_en_mem4;
  assign Mem5_instr5_MPORT_addr = Mem5_instr5_MPORT_addr_pipe_0;
  assign Mem5_instr5_MPORT_data = Mem5[Mem5_instr5_MPORT_addr]; // @[BuildingBlockNew.scala 37:25]
  assign Mem5_MPORT_4_data = io_wr_instr_mem5;
  assign Mem5_MPORT_4_addr = io_wr_en_mem5 ? wrAddr5 : PC5;
  assign Mem5_MPORT_4_mask = 1'h1;
  assign Mem5_MPORT_4_en = io_wr_en_mem5;
  assign Mem6_instr6_MPORT_addr = Mem6_instr6_MPORT_addr_pipe_0;
  assign Mem6_instr6_MPORT_data = Mem6[Mem6_instr6_MPORT_addr]; // @[BuildingBlockNew.scala 38:25]
  assign Mem6_MPORT_5_data = io_wr_instr_mem6;
  assign Mem6_MPORT_5_addr = io_wr_en_mem6 ? wrAddr6 : PC6;
  assign Mem6_MPORT_5_mask = 1'h1;
  assign Mem6_MPORT_5_en = io_wr_en_mem6;
  assign io_d_out_0_a = egress2_io_out64_0; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_0_valid_a = egress2_io_validout64_0; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_0_b = egress2_io_out64_1; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_0_valid_b = egress2_io_validout64_1; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_1_a = egress2_io_out64_2; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_1_valid_a = egress2_io_validout64_2; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_1_b = egress2_io_out64_3; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_1_valid_b = egress2_io_validout64_3; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_2_a = egress2_io_out64_4; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_2_valid_a = egress2_io_validout64_4; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_2_b = egress2_io_out64_5; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_2_valid_b = egress2_io_validout64_5; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_3_a = egress2_io_out64_6; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_3_valid_a = egress2_io_validout64_6; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_3_b = egress2_io_out64_7; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_3_valid_b = egress2_io_validout64_7; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_4_a = egress2_io_out64_8; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_4_valid_a = egress2_io_validout64_8; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_4_b = egress2_io_out64_9; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_4_valid_b = egress2_io_validout64_9; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_5_a = egress2_io_out64_10; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_5_valid_a = egress2_io_validout64_10; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_5_b = egress2_io_out64_11; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_5_valid_b = egress2_io_validout64_11; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_6_a = egress2_io_out64_12; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_6_valid_a = egress2_io_validout64_12; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_6_b = egress2_io_out64_13; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_6_valid_b = egress2_io_validout64_13; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_7_a = egress2_io_out64_14; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_7_valid_a = egress2_io_validout64_14; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_7_b = egress2_io_out64_15; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_7_valid_b = egress2_io_validout64_15; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_8_a = egress2_io_out64_16; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_8_valid_a = egress2_io_validout64_16; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_8_b = egress2_io_out64_17; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_8_valid_b = egress2_io_validout64_17; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_9_a = egress2_io_out64_18; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_9_valid_a = egress2_io_validout64_18; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_9_b = egress2_io_out64_19; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_9_valid_b = egress2_io_validout64_19; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_10_a = egress2_io_out64_20; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_10_valid_a = egress2_io_validout64_20; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_10_b = egress2_io_out64_21; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_10_valid_b = egress2_io_validout64_21; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_11_a = egress2_io_out64_22; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_11_valid_a = egress2_io_validout64_22; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_11_b = egress2_io_out64_23; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_11_valid_b = egress2_io_validout64_23; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_12_a = egress2_io_out64_24; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_12_valid_a = egress2_io_validout64_24; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_12_b = egress2_io_out64_25; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_12_valid_b = egress2_io_validout64_25; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_13_a = egress2_io_out64_26; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_13_valid_a = egress2_io_validout64_26; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_13_b = egress2_io_out64_27; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_13_valid_b = egress2_io_validout64_27; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_14_a = egress2_io_out64_28; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_14_valid_a = egress2_io_validout64_28; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_14_b = egress2_io_out64_29; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_14_valid_b = egress2_io_validout64_29; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_15_a = egress2_io_out64_30; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_15_valid_a = egress2_io_validout64_30; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_15_b = egress2_io_out64_31; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_15_valid_b = egress2_io_validout64_31; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_16_a = egress2_io_out64_32; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_16_valid_a = egress2_io_validout64_32; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_16_b = egress2_io_out64_33; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_16_valid_b = egress2_io_validout64_33; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_17_a = egress2_io_out64_34; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_17_valid_a = egress2_io_validout64_34; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_17_b = egress2_io_out64_35; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_17_valid_b = egress2_io_validout64_35; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_18_a = egress2_io_out64_36; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_18_valid_a = egress2_io_validout64_36; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_18_b = egress2_io_out64_37; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_18_valid_b = egress2_io_validout64_37; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_19_a = egress2_io_out64_38; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_19_valid_a = egress2_io_validout64_38; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_19_b = egress2_io_out64_39; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_19_valid_b = egress2_io_validout64_39; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_20_a = egress2_io_out64_40; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_20_valid_a = egress2_io_validout64_40; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_20_b = egress2_io_out64_41; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_20_valid_b = egress2_io_validout64_41; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_21_a = egress2_io_out64_42; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_21_valid_a = egress2_io_validout64_42; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_21_b = egress2_io_out64_43; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_21_valid_b = egress2_io_validout64_43; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_22_a = egress2_io_out64_44; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_22_valid_a = egress2_io_validout64_44; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_22_b = egress2_io_out64_45; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_22_valid_b = egress2_io_validout64_45; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_23_a = egress2_io_out64_46; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_23_valid_a = egress2_io_validout64_46; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_23_b = egress2_io_out64_47; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_23_valid_b = egress2_io_validout64_47; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_24_a = egress2_io_out64_48; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_24_valid_a = egress2_io_validout64_48; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_24_b = egress2_io_out64_49; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_24_valid_b = egress2_io_validout64_49; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_25_a = egress2_io_out64_50; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_25_valid_a = egress2_io_validout64_50; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_25_b = egress2_io_out64_51; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_25_valid_b = egress2_io_validout64_51; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_26_a = egress2_io_out64_52; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_26_valid_a = egress2_io_validout64_52; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_26_b = egress2_io_out64_53; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_26_valid_b = egress2_io_validout64_53; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_27_a = egress2_io_out64_54; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_27_valid_a = egress2_io_validout64_54; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_27_b = egress2_io_out64_55; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_27_valid_b = egress2_io_validout64_55; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_28_a = egress2_io_out64_56; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_28_valid_a = egress2_io_validout64_56; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_28_b = egress2_io_out64_57; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_28_valid_b = egress2_io_validout64_57; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_29_a = egress2_io_out64_58; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_29_valid_a = egress2_io_validout64_58; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_29_b = egress2_io_out64_59; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_29_valid_b = egress2_io_validout64_59; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_30_a = egress2_io_out64_60; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_30_valid_a = egress2_io_validout64_60; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_30_b = egress2_io_out64_61; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_30_valid_b = egress2_io_validout64_61; // @[BuildingBlockNew.scala 316:25]
  assign io_d_out_31_a = egress2_io_out64_62; // @[BuildingBlockNew.scala 313:19]
  assign io_d_out_31_valid_a = egress2_io_validout64_62; // @[BuildingBlockNew.scala 315:25]
  assign io_d_out_31_b = egress2_io_out64_63; // @[BuildingBlockNew.scala 314:19]
  assign io_d_out_31_valid_b = egress2_io_validout64_63; // @[BuildingBlockNew.scala 316:25]
  assign io_PC6_out = PC6; // @[BuildingBlockNew.scala 161:14]
  assign io_Addr_out = egress2_io_addrout; // @[BuildingBlockNew.scala 319:15]
  assign peCol_clock = clock;
  assign peCol_reset = reset;
  assign peCol_io_d_in_0_a = io_d_in_0_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_0_valid_a = io_d_in_0_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_0_b = io_d_in_0_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_0_valid_b = io_d_in_0_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_1_a = io_d_in_1_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_1_valid_a = io_d_in_1_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_1_b = io_d_in_1_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_1_valid_b = io_d_in_1_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_2_a = io_d_in_2_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_2_valid_a = io_d_in_2_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_2_b = io_d_in_2_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_2_valid_b = io_d_in_2_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_3_a = io_d_in_3_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_3_valid_a = io_d_in_3_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_3_b = io_d_in_3_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_3_valid_b = io_d_in_3_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_4_a = io_d_in_4_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_4_valid_a = io_d_in_4_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_4_b = io_d_in_4_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_4_valid_b = io_d_in_4_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_5_a = io_d_in_5_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_5_valid_a = io_d_in_5_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_5_b = io_d_in_5_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_5_valid_b = io_d_in_5_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_6_a = io_d_in_6_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_6_valid_a = io_d_in_6_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_6_b = io_d_in_6_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_6_valid_b = io_d_in_6_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_7_a = io_d_in_7_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_7_valid_a = io_d_in_7_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_7_b = io_d_in_7_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_7_valid_b = io_d_in_7_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_8_a = io_d_in_8_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_8_valid_a = io_d_in_8_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_8_b = io_d_in_8_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_8_valid_b = io_d_in_8_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_9_a = io_d_in_9_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_9_valid_a = io_d_in_9_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_9_b = io_d_in_9_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_9_valid_b = io_d_in_9_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_10_a = io_d_in_10_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_10_valid_a = io_d_in_10_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_10_b = io_d_in_10_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_10_valid_b = io_d_in_10_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_11_a = io_d_in_11_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_11_valid_a = io_d_in_11_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_11_b = io_d_in_11_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_11_valid_b = io_d_in_11_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_12_a = io_d_in_12_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_12_valid_a = io_d_in_12_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_12_b = io_d_in_12_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_12_valid_b = io_d_in_12_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_13_a = io_d_in_13_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_13_valid_a = io_d_in_13_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_13_b = io_d_in_13_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_13_valid_b = io_d_in_13_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_14_a = io_d_in_14_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_14_valid_a = io_d_in_14_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_14_b = io_d_in_14_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_14_valid_b = io_d_in_14_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_15_a = io_d_in_15_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_15_valid_a = io_d_in_15_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_15_b = io_d_in_15_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_15_valid_b = io_d_in_15_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_16_a = io_d_in_16_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_16_valid_a = io_d_in_16_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_16_b = io_d_in_16_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_16_valid_b = io_d_in_16_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_17_a = io_d_in_17_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_17_valid_a = io_d_in_17_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_17_b = io_d_in_17_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_17_valid_b = io_d_in_17_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_18_a = io_d_in_18_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_18_valid_a = io_d_in_18_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_18_b = io_d_in_18_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_18_valid_b = io_d_in_18_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_19_a = io_d_in_19_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_19_valid_a = io_d_in_19_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_19_b = io_d_in_19_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_19_valid_b = io_d_in_19_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_20_a = io_d_in_20_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_20_valid_a = io_d_in_20_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_20_b = io_d_in_20_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_20_valid_b = io_d_in_20_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_21_a = io_d_in_21_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_21_valid_a = io_d_in_21_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_21_b = io_d_in_21_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_21_valid_b = io_d_in_21_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_22_a = io_d_in_22_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_22_valid_a = io_d_in_22_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_22_b = io_d_in_22_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_22_valid_b = io_d_in_22_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_23_a = io_d_in_23_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_23_valid_a = io_d_in_23_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_23_b = io_d_in_23_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_23_valid_b = io_d_in_23_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_24_a = io_d_in_24_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_24_valid_a = io_d_in_24_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_24_b = io_d_in_24_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_24_valid_b = io_d_in_24_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_25_a = io_d_in_25_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_25_valid_a = io_d_in_25_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_25_b = io_d_in_25_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_25_valid_b = io_d_in_25_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_26_a = io_d_in_26_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_26_valid_a = io_d_in_26_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_26_b = io_d_in_26_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_26_valid_b = io_d_in_26_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_27_a = io_d_in_27_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_27_valid_a = io_d_in_27_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_27_b = io_d_in_27_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_27_valid_b = io_d_in_27_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_28_a = io_d_in_28_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_28_valid_a = io_d_in_28_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_28_b = io_d_in_28_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_28_valid_b = io_d_in_28_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_29_a = io_d_in_29_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_29_valid_a = io_d_in_29_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_29_b = io_d_in_29_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_29_valid_b = io_d_in_29_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_30_a = io_d_in_30_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_30_valid_a = io_d_in_30_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_30_b = io_d_in_30_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_30_valid_b = io_d_in_30_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_31_a = io_d_in_31_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_31_valid_a = io_d_in_31_valid_a; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_31_b = io_d_in_31_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_d_in_31_valid_b = io_d_in_31_valid_b; // @[BuildingBlockNew.scala 280:17]
  assign peCol_io_addrin = io_Addr_in; // @[BuildingBlockNew.scala 282:19]
  assign peCol_io_instr = Mem1_instr1_MPORT_data; // @[BuildingBlockNew.scala 223:22 BuildingBlockNew.scala 229:12]
  assign ingress1_clock = clock;
  assign ingress1_io_in64_0 = peCol_io_d_out_0_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_1 = peCol_io_d_out_0_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_2 = peCol_io_d_out_1_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_3 = peCol_io_d_out_1_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_4 = peCol_io_d_out_2_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_5 = peCol_io_d_out_2_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_6 = peCol_io_d_out_3_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_7 = peCol_io_d_out_3_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_8 = peCol_io_d_out_4_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_9 = peCol_io_d_out_4_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_10 = peCol_io_d_out_5_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_11 = peCol_io_d_out_5_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_12 = peCol_io_d_out_6_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_13 = peCol_io_d_out_6_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_14 = peCol_io_d_out_7_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_15 = peCol_io_d_out_7_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_16 = peCol_io_d_out_8_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_17 = peCol_io_d_out_8_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_18 = peCol_io_d_out_9_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_19 = peCol_io_d_out_9_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_20 = peCol_io_d_out_10_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_21 = peCol_io_d_out_10_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_22 = peCol_io_d_out_11_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_23 = peCol_io_d_out_11_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_24 = peCol_io_d_out_12_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_25 = peCol_io_d_out_12_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_26 = peCol_io_d_out_13_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_27 = peCol_io_d_out_13_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_28 = peCol_io_d_out_14_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_29 = peCol_io_d_out_14_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_30 = peCol_io_d_out_15_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_31 = peCol_io_d_out_15_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_32 = peCol_io_d_out_16_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_33 = peCol_io_d_out_16_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_34 = peCol_io_d_out_17_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_35 = peCol_io_d_out_17_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_36 = peCol_io_d_out_18_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_37 = peCol_io_d_out_18_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_38 = peCol_io_d_out_19_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_39 = peCol_io_d_out_19_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_40 = peCol_io_d_out_20_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_41 = peCol_io_d_out_20_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_42 = peCol_io_d_out_21_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_43 = peCol_io_d_out_21_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_44 = peCol_io_d_out_22_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_45 = peCol_io_d_out_22_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_46 = peCol_io_d_out_23_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_47 = peCol_io_d_out_23_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_48 = peCol_io_d_out_24_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_49 = peCol_io_d_out_24_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_50 = peCol_io_d_out_25_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_51 = peCol_io_d_out_25_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_52 = peCol_io_d_out_26_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_53 = peCol_io_d_out_26_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_54 = peCol_io_d_out_27_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_55 = peCol_io_d_out_27_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_56 = peCol_io_d_out_28_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_57 = peCol_io_d_out_28_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_58 = peCol_io_d_out_29_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_59 = peCol_io_d_out_29_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_60 = peCol_io_d_out_30_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_61 = peCol_io_d_out_30_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_in64_62 = peCol_io_d_out_31_a; // @[BuildingBlockNew.scala 287:27]
  assign ingress1_io_in64_63 = peCol_io_d_out_31_b; // @[BuildingBlockNew.scala 288:29]
  assign ingress1_io_validin64_0 = peCol_io_d_out_0_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_1 = peCol_io_d_out_0_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_2 = peCol_io_d_out_1_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_3 = peCol_io_d_out_1_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_4 = peCol_io_d_out_2_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_5 = peCol_io_d_out_2_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_6 = peCol_io_d_out_3_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_7 = peCol_io_d_out_3_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_8 = peCol_io_d_out_4_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_9 = peCol_io_d_out_4_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_10 = peCol_io_d_out_5_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_11 = peCol_io_d_out_5_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_12 = peCol_io_d_out_6_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_13 = peCol_io_d_out_6_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_14 = peCol_io_d_out_7_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_15 = peCol_io_d_out_7_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_16 = peCol_io_d_out_8_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_17 = peCol_io_d_out_8_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_18 = peCol_io_d_out_9_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_19 = peCol_io_d_out_9_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_20 = peCol_io_d_out_10_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_21 = peCol_io_d_out_10_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_22 = peCol_io_d_out_11_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_23 = peCol_io_d_out_11_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_24 = peCol_io_d_out_12_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_25 = peCol_io_d_out_12_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_26 = peCol_io_d_out_13_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_27 = peCol_io_d_out_13_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_28 = peCol_io_d_out_14_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_29 = peCol_io_d_out_14_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_30 = peCol_io_d_out_15_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_31 = peCol_io_d_out_15_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_32 = peCol_io_d_out_16_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_33 = peCol_io_d_out_16_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_34 = peCol_io_d_out_17_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_35 = peCol_io_d_out_17_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_36 = peCol_io_d_out_18_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_37 = peCol_io_d_out_18_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_38 = peCol_io_d_out_19_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_39 = peCol_io_d_out_19_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_40 = peCol_io_d_out_20_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_41 = peCol_io_d_out_20_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_42 = peCol_io_d_out_21_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_43 = peCol_io_d_out_21_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_44 = peCol_io_d_out_22_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_45 = peCol_io_d_out_22_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_46 = peCol_io_d_out_23_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_47 = peCol_io_d_out_23_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_48 = peCol_io_d_out_24_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_49 = peCol_io_d_out_24_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_50 = peCol_io_d_out_25_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_51 = peCol_io_d_out_25_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_52 = peCol_io_d_out_26_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_53 = peCol_io_d_out_26_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_54 = peCol_io_d_out_27_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_55 = peCol_io_d_out_27_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_56 = peCol_io_d_out_28_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_57 = peCol_io_d_out_28_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_58 = peCol_io_d_out_29_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_59 = peCol_io_d_out_29_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_60 = peCol_io_d_out_30_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_61 = peCol_io_d_out_30_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_validin64_62 = peCol_io_d_out_31_valid_a; // @[BuildingBlockNew.scala 289:32]
  assign ingress1_io_validin64_63 = peCol_io_d_out_31_valid_b; // @[BuildingBlockNew.scala 290:34]
  assign ingress1_io_addrin = peCol_io_addrout; // @[BuildingBlockNew.scala 285:22]
  assign ingress1_io_ctrl = Mem2_instr2_MPORT_data; // @[BuildingBlockNew.scala 232:22 BuildingBlockNew.scala 238:12]
  assign ingress2_clock = clock;
  assign ingress2_io_in64_0 = ingress1_io_out64_0; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_1 = ingress1_io_out64_1; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_2 = ingress1_io_out64_2; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_3 = ingress1_io_out64_3; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_4 = ingress1_io_out64_4; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_5 = ingress1_io_out64_5; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_6 = ingress1_io_out64_6; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_7 = ingress1_io_out64_7; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_8 = ingress1_io_out64_8; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_9 = ingress1_io_out64_9; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_10 = ingress1_io_out64_10; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_11 = ingress1_io_out64_11; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_12 = ingress1_io_out64_12; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_13 = ingress1_io_out64_13; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_14 = ingress1_io_out64_14; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_15 = ingress1_io_out64_15; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_16 = ingress1_io_out64_16; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_17 = ingress1_io_out64_17; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_18 = ingress1_io_out64_18; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_19 = ingress1_io_out64_19; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_20 = ingress1_io_out64_20; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_21 = ingress1_io_out64_21; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_22 = ingress1_io_out64_22; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_23 = ingress1_io_out64_23; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_24 = ingress1_io_out64_24; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_25 = ingress1_io_out64_25; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_26 = ingress1_io_out64_26; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_27 = ingress1_io_out64_27; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_28 = ingress1_io_out64_28; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_29 = ingress1_io_out64_29; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_30 = ingress1_io_out64_30; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_31 = ingress1_io_out64_31; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_32 = ingress1_io_out64_32; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_33 = ingress1_io_out64_33; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_34 = ingress1_io_out64_34; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_35 = ingress1_io_out64_35; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_36 = ingress1_io_out64_36; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_37 = ingress1_io_out64_37; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_38 = ingress1_io_out64_38; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_39 = ingress1_io_out64_39; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_40 = ingress1_io_out64_40; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_41 = ingress1_io_out64_41; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_42 = ingress1_io_out64_42; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_43 = ingress1_io_out64_43; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_44 = ingress1_io_out64_44; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_45 = ingress1_io_out64_45; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_46 = ingress1_io_out64_46; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_47 = ingress1_io_out64_47; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_48 = ingress1_io_out64_48; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_49 = ingress1_io_out64_49; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_50 = ingress1_io_out64_50; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_51 = ingress1_io_out64_51; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_52 = ingress1_io_out64_52; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_53 = ingress1_io_out64_53; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_54 = ingress1_io_out64_54; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_55 = ingress1_io_out64_55; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_56 = ingress1_io_out64_56; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_57 = ingress1_io_out64_57; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_58 = ingress1_io_out64_58; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_59 = ingress1_io_out64_59; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_60 = ingress1_io_out64_60; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_61 = ingress1_io_out64_61; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_62 = ingress1_io_out64_62; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_in64_63 = ingress1_io_out64_63; // @[BuildingBlockNew.scala 293:20]
  assign ingress2_io_validin64_0 = ingress1_io_validout64_0; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_1 = ingress1_io_validout64_1; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_2 = ingress1_io_validout64_2; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_3 = ingress1_io_validout64_3; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_4 = ingress1_io_validout64_4; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_5 = ingress1_io_validout64_5; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_6 = ingress1_io_validout64_6; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_7 = ingress1_io_validout64_7; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_8 = ingress1_io_validout64_8; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_9 = ingress1_io_validout64_9; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_10 = ingress1_io_validout64_10; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_11 = ingress1_io_validout64_11; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_12 = ingress1_io_validout64_12; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_13 = ingress1_io_validout64_13; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_14 = ingress1_io_validout64_14; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_15 = ingress1_io_validout64_15; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_16 = ingress1_io_validout64_16; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_17 = ingress1_io_validout64_17; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_18 = ingress1_io_validout64_18; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_19 = ingress1_io_validout64_19; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_20 = ingress1_io_validout64_20; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_21 = ingress1_io_validout64_21; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_22 = ingress1_io_validout64_22; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_23 = ingress1_io_validout64_23; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_24 = ingress1_io_validout64_24; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_25 = ingress1_io_validout64_25; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_26 = ingress1_io_validout64_26; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_27 = ingress1_io_validout64_27; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_28 = ingress1_io_validout64_28; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_29 = ingress1_io_validout64_29; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_30 = ingress1_io_validout64_30; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_31 = ingress1_io_validout64_31; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_32 = ingress1_io_validout64_32; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_33 = ingress1_io_validout64_33; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_34 = ingress1_io_validout64_34; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_35 = ingress1_io_validout64_35; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_36 = ingress1_io_validout64_36; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_37 = ingress1_io_validout64_37; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_38 = ingress1_io_validout64_38; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_39 = ingress1_io_validout64_39; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_40 = ingress1_io_validout64_40; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_41 = ingress1_io_validout64_41; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_42 = ingress1_io_validout64_42; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_43 = ingress1_io_validout64_43; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_44 = ingress1_io_validout64_44; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_45 = ingress1_io_validout64_45; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_46 = ingress1_io_validout64_46; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_47 = ingress1_io_validout64_47; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_48 = ingress1_io_validout64_48; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_49 = ingress1_io_validout64_49; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_50 = ingress1_io_validout64_50; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_51 = ingress1_io_validout64_51; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_52 = ingress1_io_validout64_52; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_53 = ingress1_io_validout64_53; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_54 = ingress1_io_validout64_54; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_55 = ingress1_io_validout64_55; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_56 = ingress1_io_validout64_56; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_57 = ingress1_io_validout64_57; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_58 = ingress1_io_validout64_58; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_59 = ingress1_io_validout64_59; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_60 = ingress1_io_validout64_60; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_61 = ingress1_io_validout64_61; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_62 = ingress1_io_validout64_62; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_validin64_63 = ingress1_io_validout64_63; // @[BuildingBlockNew.scala 294:25]
  assign ingress2_io_addrin = ingress1_io_addrout; // @[BuildingBlockNew.scala 296:22]
  assign ingress2_io_ctrl = Mem3_instr3_MPORT_data; // @[BuildingBlockNew.scala 241:22 BuildingBlockNew.scala 247:12]
  assign middle_clock = clock;
  assign middle_io_in64_0 = ingress2_io_out64_0; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_1 = ingress2_io_out64_1; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_2 = ingress2_io_out64_2; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_3 = ingress2_io_out64_3; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_4 = ingress2_io_out64_4; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_5 = ingress2_io_out64_5; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_6 = ingress2_io_out64_6; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_7 = ingress2_io_out64_7; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_8 = ingress2_io_out64_8; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_9 = ingress2_io_out64_9; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_10 = ingress2_io_out64_10; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_11 = ingress2_io_out64_11; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_12 = ingress2_io_out64_12; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_13 = ingress2_io_out64_13; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_14 = ingress2_io_out64_14; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_15 = ingress2_io_out64_15; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_16 = ingress2_io_out64_16; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_17 = ingress2_io_out64_17; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_18 = ingress2_io_out64_18; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_19 = ingress2_io_out64_19; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_20 = ingress2_io_out64_20; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_21 = ingress2_io_out64_21; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_22 = ingress2_io_out64_22; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_23 = ingress2_io_out64_23; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_24 = ingress2_io_out64_24; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_25 = ingress2_io_out64_25; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_26 = ingress2_io_out64_26; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_27 = ingress2_io_out64_27; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_28 = ingress2_io_out64_28; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_29 = ingress2_io_out64_29; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_30 = ingress2_io_out64_30; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_31 = ingress2_io_out64_31; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_32 = ingress2_io_out64_32; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_33 = ingress2_io_out64_33; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_34 = ingress2_io_out64_34; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_35 = ingress2_io_out64_35; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_36 = ingress2_io_out64_36; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_37 = ingress2_io_out64_37; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_38 = ingress2_io_out64_38; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_39 = ingress2_io_out64_39; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_40 = ingress2_io_out64_40; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_41 = ingress2_io_out64_41; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_42 = ingress2_io_out64_42; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_43 = ingress2_io_out64_43; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_44 = ingress2_io_out64_44; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_45 = ingress2_io_out64_45; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_46 = ingress2_io_out64_46; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_47 = ingress2_io_out64_47; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_48 = ingress2_io_out64_48; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_49 = ingress2_io_out64_49; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_50 = ingress2_io_out64_50; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_51 = ingress2_io_out64_51; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_52 = ingress2_io_out64_52; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_53 = ingress2_io_out64_53; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_54 = ingress2_io_out64_54; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_55 = ingress2_io_out64_55; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_56 = ingress2_io_out64_56; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_57 = ingress2_io_out64_57; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_58 = ingress2_io_out64_58; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_59 = ingress2_io_out64_59; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_60 = ingress2_io_out64_60; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_61 = ingress2_io_out64_61; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_62 = ingress2_io_out64_62; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_in64_63 = ingress2_io_out64_63; // @[BuildingBlockNew.scala 297:18]
  assign middle_io_validin64_0 = ingress2_io_validout64_0; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_1 = ingress2_io_validout64_1; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_2 = ingress2_io_validout64_2; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_3 = ingress2_io_validout64_3; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_4 = ingress2_io_validout64_4; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_5 = ingress2_io_validout64_5; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_6 = ingress2_io_validout64_6; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_7 = ingress2_io_validout64_7; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_8 = ingress2_io_validout64_8; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_9 = ingress2_io_validout64_9; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_10 = ingress2_io_validout64_10; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_11 = ingress2_io_validout64_11; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_12 = ingress2_io_validout64_12; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_13 = ingress2_io_validout64_13; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_14 = ingress2_io_validout64_14; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_15 = ingress2_io_validout64_15; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_16 = ingress2_io_validout64_16; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_17 = ingress2_io_validout64_17; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_18 = ingress2_io_validout64_18; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_19 = ingress2_io_validout64_19; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_20 = ingress2_io_validout64_20; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_21 = ingress2_io_validout64_21; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_22 = ingress2_io_validout64_22; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_23 = ingress2_io_validout64_23; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_24 = ingress2_io_validout64_24; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_25 = ingress2_io_validout64_25; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_26 = ingress2_io_validout64_26; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_27 = ingress2_io_validout64_27; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_28 = ingress2_io_validout64_28; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_29 = ingress2_io_validout64_29; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_30 = ingress2_io_validout64_30; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_31 = ingress2_io_validout64_31; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_32 = ingress2_io_validout64_32; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_33 = ingress2_io_validout64_33; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_34 = ingress2_io_validout64_34; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_35 = ingress2_io_validout64_35; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_36 = ingress2_io_validout64_36; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_37 = ingress2_io_validout64_37; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_38 = ingress2_io_validout64_38; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_39 = ingress2_io_validout64_39; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_40 = ingress2_io_validout64_40; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_41 = ingress2_io_validout64_41; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_42 = ingress2_io_validout64_42; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_43 = ingress2_io_validout64_43; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_44 = ingress2_io_validout64_44; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_45 = ingress2_io_validout64_45; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_46 = ingress2_io_validout64_46; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_47 = ingress2_io_validout64_47; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_48 = ingress2_io_validout64_48; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_49 = ingress2_io_validout64_49; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_50 = ingress2_io_validout64_50; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_51 = ingress2_io_validout64_51; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_52 = ingress2_io_validout64_52; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_53 = ingress2_io_validout64_53; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_54 = ingress2_io_validout64_54; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_55 = ingress2_io_validout64_55; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_56 = ingress2_io_validout64_56; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_57 = ingress2_io_validout64_57; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_58 = ingress2_io_validout64_58; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_59 = ingress2_io_validout64_59; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_60 = ingress2_io_validout64_60; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_61 = ingress2_io_validout64_61; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_62 = ingress2_io_validout64_62; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_validin64_63 = ingress2_io_validout64_63; // @[BuildingBlockNew.scala 298:23]
  assign middle_io_addrin = ingress2_io_addrout; // @[BuildingBlockNew.scala 300:20]
  assign middle_io_ctrl = Mem4_instr4_MPORT_data; // @[BuildingBlockNew.scala 250:22 BuildingBlockNew.scala 256:12]
  assign egress1_clock = clock;
  assign egress1_io_in64_0 = middle_io_out64_0; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_1 = middle_io_out64_1; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_2 = middle_io_out64_2; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_3 = middle_io_out64_3; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_4 = middle_io_out64_4; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_5 = middle_io_out64_5; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_6 = middle_io_out64_6; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_7 = middle_io_out64_7; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_8 = middle_io_out64_8; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_9 = middle_io_out64_9; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_10 = middle_io_out64_10; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_11 = middle_io_out64_11; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_12 = middle_io_out64_12; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_13 = middle_io_out64_13; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_14 = middle_io_out64_14; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_15 = middle_io_out64_15; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_16 = middle_io_out64_16; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_17 = middle_io_out64_17; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_18 = middle_io_out64_18; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_19 = middle_io_out64_19; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_20 = middle_io_out64_20; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_21 = middle_io_out64_21; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_22 = middle_io_out64_22; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_23 = middle_io_out64_23; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_24 = middle_io_out64_24; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_25 = middle_io_out64_25; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_26 = middle_io_out64_26; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_27 = middle_io_out64_27; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_28 = middle_io_out64_28; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_29 = middle_io_out64_29; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_30 = middle_io_out64_30; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_31 = middle_io_out64_31; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_32 = middle_io_out64_32; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_33 = middle_io_out64_33; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_34 = middle_io_out64_34; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_35 = middle_io_out64_35; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_36 = middle_io_out64_36; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_37 = middle_io_out64_37; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_38 = middle_io_out64_38; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_39 = middle_io_out64_39; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_40 = middle_io_out64_40; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_41 = middle_io_out64_41; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_42 = middle_io_out64_42; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_43 = middle_io_out64_43; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_44 = middle_io_out64_44; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_45 = middle_io_out64_45; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_46 = middle_io_out64_46; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_47 = middle_io_out64_47; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_48 = middle_io_out64_48; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_49 = middle_io_out64_49; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_50 = middle_io_out64_50; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_51 = middle_io_out64_51; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_52 = middle_io_out64_52; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_53 = middle_io_out64_53; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_54 = middle_io_out64_54; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_55 = middle_io_out64_55; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_56 = middle_io_out64_56; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_57 = middle_io_out64_57; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_58 = middle_io_out64_58; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_59 = middle_io_out64_59; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_60 = middle_io_out64_60; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_61 = middle_io_out64_61; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_62 = middle_io_out64_62; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_in64_63 = middle_io_out64_63; // @[BuildingBlockNew.scala 301:19]
  assign egress1_io_validin64_0 = middle_io_validout64_0; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_1 = middle_io_validout64_1; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_2 = middle_io_validout64_2; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_3 = middle_io_validout64_3; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_4 = middle_io_validout64_4; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_5 = middle_io_validout64_5; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_6 = middle_io_validout64_6; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_7 = middle_io_validout64_7; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_8 = middle_io_validout64_8; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_9 = middle_io_validout64_9; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_10 = middle_io_validout64_10; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_11 = middle_io_validout64_11; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_12 = middle_io_validout64_12; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_13 = middle_io_validout64_13; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_14 = middle_io_validout64_14; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_15 = middle_io_validout64_15; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_16 = middle_io_validout64_16; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_17 = middle_io_validout64_17; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_18 = middle_io_validout64_18; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_19 = middle_io_validout64_19; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_20 = middle_io_validout64_20; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_21 = middle_io_validout64_21; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_22 = middle_io_validout64_22; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_23 = middle_io_validout64_23; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_24 = middle_io_validout64_24; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_25 = middle_io_validout64_25; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_26 = middle_io_validout64_26; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_27 = middle_io_validout64_27; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_28 = middle_io_validout64_28; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_29 = middle_io_validout64_29; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_30 = middle_io_validout64_30; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_31 = middle_io_validout64_31; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_32 = middle_io_validout64_32; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_33 = middle_io_validout64_33; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_34 = middle_io_validout64_34; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_35 = middle_io_validout64_35; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_36 = middle_io_validout64_36; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_37 = middle_io_validout64_37; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_38 = middle_io_validout64_38; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_39 = middle_io_validout64_39; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_40 = middle_io_validout64_40; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_41 = middle_io_validout64_41; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_42 = middle_io_validout64_42; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_43 = middle_io_validout64_43; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_44 = middle_io_validout64_44; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_45 = middle_io_validout64_45; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_46 = middle_io_validout64_46; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_47 = middle_io_validout64_47; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_48 = middle_io_validout64_48; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_49 = middle_io_validout64_49; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_50 = middle_io_validout64_50; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_51 = middle_io_validout64_51; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_52 = middle_io_validout64_52; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_53 = middle_io_validout64_53; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_54 = middle_io_validout64_54; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_55 = middle_io_validout64_55; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_56 = middle_io_validout64_56; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_57 = middle_io_validout64_57; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_58 = middle_io_validout64_58; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_59 = middle_io_validout64_59; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_60 = middle_io_validout64_60; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_61 = middle_io_validout64_61; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_62 = middle_io_validout64_62; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_validin64_63 = middle_io_validout64_63; // @[BuildingBlockNew.scala 302:24]
  assign egress1_io_addrin = middle_io_addrout; // @[BuildingBlockNew.scala 304:21]
  assign egress1_io_ctrl = Mem5_instr5_MPORT_data; // @[BuildingBlockNew.scala 259:22 BuildingBlockNew.scala 265:12]
  assign egress2_clock = clock;
  assign egress2_io_in64_0 = egress1_io_out64_0; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_1 = egress1_io_out64_1; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_2 = egress1_io_out64_2; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_3 = egress1_io_out64_3; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_4 = egress1_io_out64_4; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_5 = egress1_io_out64_5; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_6 = egress1_io_out64_6; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_7 = egress1_io_out64_7; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_8 = egress1_io_out64_8; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_9 = egress1_io_out64_9; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_10 = egress1_io_out64_10; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_11 = egress1_io_out64_11; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_12 = egress1_io_out64_12; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_13 = egress1_io_out64_13; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_14 = egress1_io_out64_14; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_15 = egress1_io_out64_15; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_16 = egress1_io_out64_16; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_17 = egress1_io_out64_17; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_18 = egress1_io_out64_18; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_19 = egress1_io_out64_19; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_20 = egress1_io_out64_20; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_21 = egress1_io_out64_21; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_22 = egress1_io_out64_22; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_23 = egress1_io_out64_23; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_24 = egress1_io_out64_24; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_25 = egress1_io_out64_25; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_26 = egress1_io_out64_26; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_27 = egress1_io_out64_27; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_28 = egress1_io_out64_28; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_29 = egress1_io_out64_29; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_30 = egress1_io_out64_30; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_31 = egress1_io_out64_31; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_32 = egress1_io_out64_32; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_33 = egress1_io_out64_33; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_34 = egress1_io_out64_34; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_35 = egress1_io_out64_35; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_36 = egress1_io_out64_36; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_37 = egress1_io_out64_37; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_38 = egress1_io_out64_38; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_39 = egress1_io_out64_39; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_40 = egress1_io_out64_40; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_41 = egress1_io_out64_41; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_42 = egress1_io_out64_42; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_43 = egress1_io_out64_43; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_44 = egress1_io_out64_44; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_45 = egress1_io_out64_45; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_46 = egress1_io_out64_46; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_47 = egress1_io_out64_47; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_48 = egress1_io_out64_48; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_49 = egress1_io_out64_49; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_50 = egress1_io_out64_50; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_51 = egress1_io_out64_51; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_52 = egress1_io_out64_52; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_53 = egress1_io_out64_53; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_54 = egress1_io_out64_54; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_55 = egress1_io_out64_55; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_56 = egress1_io_out64_56; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_57 = egress1_io_out64_57; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_58 = egress1_io_out64_58; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_59 = egress1_io_out64_59; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_60 = egress1_io_out64_60; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_61 = egress1_io_out64_61; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_62 = egress1_io_out64_62; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_in64_63 = egress1_io_out64_63; // @[BuildingBlockNew.scala 305:19]
  assign egress2_io_validin64_0 = egress1_io_validout64_0; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_1 = egress1_io_validout64_1; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_2 = egress1_io_validout64_2; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_3 = egress1_io_validout64_3; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_4 = egress1_io_validout64_4; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_5 = egress1_io_validout64_5; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_6 = egress1_io_validout64_6; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_7 = egress1_io_validout64_7; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_8 = egress1_io_validout64_8; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_9 = egress1_io_validout64_9; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_10 = egress1_io_validout64_10; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_11 = egress1_io_validout64_11; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_12 = egress1_io_validout64_12; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_13 = egress1_io_validout64_13; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_14 = egress1_io_validout64_14; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_15 = egress1_io_validout64_15; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_16 = egress1_io_validout64_16; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_17 = egress1_io_validout64_17; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_18 = egress1_io_validout64_18; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_19 = egress1_io_validout64_19; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_20 = egress1_io_validout64_20; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_21 = egress1_io_validout64_21; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_22 = egress1_io_validout64_22; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_23 = egress1_io_validout64_23; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_24 = egress1_io_validout64_24; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_25 = egress1_io_validout64_25; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_26 = egress1_io_validout64_26; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_27 = egress1_io_validout64_27; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_28 = egress1_io_validout64_28; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_29 = egress1_io_validout64_29; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_30 = egress1_io_validout64_30; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_31 = egress1_io_validout64_31; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_32 = egress1_io_validout64_32; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_33 = egress1_io_validout64_33; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_34 = egress1_io_validout64_34; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_35 = egress1_io_validout64_35; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_36 = egress1_io_validout64_36; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_37 = egress1_io_validout64_37; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_38 = egress1_io_validout64_38; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_39 = egress1_io_validout64_39; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_40 = egress1_io_validout64_40; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_41 = egress1_io_validout64_41; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_42 = egress1_io_validout64_42; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_43 = egress1_io_validout64_43; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_44 = egress1_io_validout64_44; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_45 = egress1_io_validout64_45; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_46 = egress1_io_validout64_46; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_47 = egress1_io_validout64_47; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_48 = egress1_io_validout64_48; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_49 = egress1_io_validout64_49; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_50 = egress1_io_validout64_50; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_51 = egress1_io_validout64_51; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_52 = egress1_io_validout64_52; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_53 = egress1_io_validout64_53; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_54 = egress1_io_validout64_54; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_55 = egress1_io_validout64_55; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_56 = egress1_io_validout64_56; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_57 = egress1_io_validout64_57; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_58 = egress1_io_validout64_58; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_59 = egress1_io_validout64_59; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_60 = egress1_io_validout64_60; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_61 = egress1_io_validout64_61; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_62 = egress1_io_validout64_62; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_validin64_63 = egress1_io_validout64_63; // @[BuildingBlockNew.scala 306:24]
  assign egress2_io_addrin = egress1_io_addrout; // @[BuildingBlockNew.scala 308:21]
  assign egress2_io_ctrl = Mem6_instr6_MPORT_data; // @[BuildingBlockNew.scala 268:22 BuildingBlockNew.scala 274:12]
  always @(posedge clock) begin
    if(Mem1_MPORT_en & Mem1_MPORT_mask) begin
      Mem1[Mem1_MPORT_addr] <= Mem1_MPORT_data; // @[BuildingBlockNew.scala 33:25]
    end
    if (io_wr_en_mem1) begin
      Mem1_instr1_MPORT_addr_pipe_0 <= wrAddr1;
    end else begin
      Mem1_instr1_MPORT_addr_pipe_0 <= PC1;
    end
    if(Mem2_MPORT_1_en & Mem2_MPORT_1_mask) begin
      Mem2[Mem2_MPORT_1_addr] <= Mem2_MPORT_1_data; // @[BuildingBlockNew.scala 34:25]
    end
    if (io_wr_en_mem2) begin
      Mem2_instr2_MPORT_addr_pipe_0 <= wrAddr2;
    end else begin
      Mem2_instr2_MPORT_addr_pipe_0 <= PC2;
    end
    if(Mem3_MPORT_2_en & Mem3_MPORT_2_mask) begin
      Mem3[Mem3_MPORT_2_addr] <= Mem3_MPORT_2_data; // @[BuildingBlockNew.scala 35:25]
    end
    if (io_wr_en_mem3) begin
      Mem3_instr3_MPORT_addr_pipe_0 <= wrAddr3;
    end else begin
      Mem3_instr3_MPORT_addr_pipe_0 <= PC3;
    end
    if(Mem4_MPORT_3_en & Mem4_MPORT_3_mask) begin
      Mem4[Mem4_MPORT_3_addr] <= Mem4_MPORT_3_data; // @[BuildingBlockNew.scala 36:25]
    end
    if (io_wr_en_mem4) begin
      Mem4_instr4_MPORT_addr_pipe_0 <= wrAddr4;
    end else begin
      Mem4_instr4_MPORT_addr_pipe_0 <= PC4;
    end
    if(Mem5_MPORT_4_en & Mem5_MPORT_4_mask) begin
      Mem5[Mem5_MPORT_4_addr] <= Mem5_MPORT_4_data; // @[BuildingBlockNew.scala 37:25]
    end
    if (io_wr_en_mem5) begin
      Mem5_instr5_MPORT_addr_pipe_0 <= wrAddr5;
    end else begin
      Mem5_instr5_MPORT_addr_pipe_0 <= PC5;
    end
    if(Mem6_MPORT_5_en & Mem6_MPORT_5_mask) begin
      Mem6[Mem6_MPORT_5_addr] <= Mem6_MPORT_5_data; // @[BuildingBlockNew.scala 38:25]
    end
    if (io_wr_en_mem6) begin
      Mem6_instr6_MPORT_addr_pipe_0 <= wrAddr6;
    end else begin
      Mem6_instr6_MPORT_addr_pipe_0 <= PC6;
    end
    if (reset) begin // @[BuildingBlockNew.scala 39:20]
      PC1 <= 8'h0; // @[BuildingBlockNew.scala 39:20]
    end else begin
      PC1 <= io_PC1_in; // @[BuildingBlockNew.scala 154:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 40:20]
      PC2 <= 8'h0; // @[BuildingBlockNew.scala 40:20]
    end else begin
      PC2 <= PC1; // @[BuildingBlockNew.scala 155:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 41:20]
      PC3 <= 8'h0; // @[BuildingBlockNew.scala 41:20]
    end else begin
      PC3 <= PC2; // @[BuildingBlockNew.scala 156:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 42:20]
      PC4 <= 8'h0; // @[BuildingBlockNew.scala 42:20]
    end else begin
      PC4 <= PC3; // @[BuildingBlockNew.scala 157:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 43:20]
      PC5 <= 8'h0; // @[BuildingBlockNew.scala 43:20]
    end else begin
      PC5 <= PC4; // @[BuildingBlockNew.scala 158:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 44:20]
      PC6 <= 8'h0; // @[BuildingBlockNew.scala 44:20]
    end else begin
      PC6 <= PC5; // @[BuildingBlockNew.scala 159:7]
    end
    if (reset) begin // @[BuildingBlockNew.scala 45:24]
      wrAddr1 <= 8'h0; // @[BuildingBlockNew.scala 45:24]
    end else if (io_wr_en_mem1) begin // @[BuildingBlockNew.scala 223:22]
      wrAddr1 <= _wrAddr1_T_1; // @[BuildingBlockNew.scala 226:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 46:24]
      wrAddr2 <= 8'h0; // @[BuildingBlockNew.scala 46:24]
    end else if (io_wr_en_mem2) begin // @[BuildingBlockNew.scala 232:22]
      wrAddr2 <= _wrAddr2_T_1; // @[BuildingBlockNew.scala 235:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 47:24]
      wrAddr3 <= 8'h0; // @[BuildingBlockNew.scala 47:24]
    end else if (io_wr_en_mem3) begin // @[BuildingBlockNew.scala 241:22]
      wrAddr3 <= _wrAddr3_T_1; // @[BuildingBlockNew.scala 244:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 48:24]
      wrAddr4 <= 8'h0; // @[BuildingBlockNew.scala 48:24]
    end else if (io_wr_en_mem4) begin // @[BuildingBlockNew.scala 250:22]
      wrAddr4 <= _wrAddr4_T_1; // @[BuildingBlockNew.scala 253:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 49:24]
      wrAddr5 <= 8'h0; // @[BuildingBlockNew.scala 49:24]
    end else if (io_wr_en_mem5) begin // @[BuildingBlockNew.scala 259:22]
      wrAddr5 <= _wrAddr5_T_1; // @[BuildingBlockNew.scala 262:13]
    end
    if (reset) begin // @[BuildingBlockNew.scala 50:24]
      wrAddr6 <= 8'h0; // @[BuildingBlockNew.scala 50:24]
    end else if (io_wr_en_mem6) begin // @[BuildingBlockNew.scala 268:22]
      wrAddr6 <= _wrAddr6_T_1; // @[BuildingBlockNew.scala 271:13]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {9{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    Mem1[initvar] = _RAND_0[287:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    Mem2[initvar] = _RAND_2[127:0];
  _RAND_4 = {4{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    Mem3[initvar] = _RAND_4[127:0];
  _RAND_6 = {4{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    Mem4[initvar] = _RAND_6[127:0];
  _RAND_8 = {4{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    Mem5[initvar] = _RAND_8[127:0];
  _RAND_10 = {4{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    Mem6[initvar] = _RAND_10[127:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  Mem1_instr1_MPORT_addr_pipe_0 = _RAND_1[7:0];
  _RAND_3 = {1{`RANDOM}};
  Mem2_instr2_MPORT_addr_pipe_0 = _RAND_3[7:0];
  _RAND_5 = {1{`RANDOM}};
  Mem3_instr3_MPORT_addr_pipe_0 = _RAND_5[7:0];
  _RAND_7 = {1{`RANDOM}};
  Mem4_instr4_MPORT_addr_pipe_0 = _RAND_7[7:0];
  _RAND_9 = {1{`RANDOM}};
  Mem5_instr5_MPORT_addr_pipe_0 = _RAND_9[7:0];
  _RAND_11 = {1{`RANDOM}};
  Mem6_instr6_MPORT_addr_pipe_0 = _RAND_11[7:0];
  _RAND_12 = {1{`RANDOM}};
  PC1 = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  PC2 = _RAND_13[7:0];
  _RAND_14 = {1{`RANDOM}};
  PC3 = _RAND_14[7:0];
  _RAND_15 = {1{`RANDOM}};
  PC4 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  PC5 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  PC6 = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  wrAddr1 = _RAND_18[7:0];
  _RAND_19 = {1{`RANDOM}};
  wrAddr2 = _RAND_19[7:0];
  _RAND_20 = {1{`RANDOM}};
  wrAddr3 = _RAND_20[7:0];
  _RAND_21 = {1{`RANDOM}};
  wrAddr4 = _RAND_21[7:0];
  _RAND_22 = {1{`RANDOM}};
  wrAddr5 = _RAND_22[7:0];
  _RAND_23 = {1{`RANDOM}};
  wrAddr6 = _RAND_23[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module BP(
  input          clock,
  input          reset,
  input          io_wr_en_mem1_0,
  input          io_wr_en_mem1_1,
  input          io_wr_en_mem1_2,
  input          io_wr_en_mem1_3,
  input          io_wr_en_mem1_4,
  input          io_wr_en_mem1_5,
  input          io_wr_en_mem1_6,
  input          io_wr_en_mem1_7,
  input          io_wr_en_mem1_8,
  input          io_wr_en_mem1_9,
  input          io_wr_en_mem1_10,
  input          io_wr_en_mem1_11,
  input          io_wr_en_mem1_12,
  input          io_wr_en_mem1_13,
  input          io_wr_en_mem1_14,
  input          io_wr_en_mem1_15,
  input          io_wr_en_mem1_16,
  input          io_wr_en_mem1_17,
  input          io_wr_en_mem1_18,
  input          io_wr_en_mem1_19,
  input          io_wr_en_mem1_20,
  input          io_wr_en_mem2_0,
  input          io_wr_en_mem2_1,
  input          io_wr_en_mem2_2,
  input          io_wr_en_mem2_3,
  input          io_wr_en_mem2_4,
  input          io_wr_en_mem2_5,
  input          io_wr_en_mem2_6,
  input          io_wr_en_mem2_7,
  input          io_wr_en_mem2_8,
  input          io_wr_en_mem2_9,
  input          io_wr_en_mem2_10,
  input          io_wr_en_mem2_11,
  input          io_wr_en_mem2_12,
  input          io_wr_en_mem2_13,
  input          io_wr_en_mem2_14,
  input          io_wr_en_mem2_15,
  input          io_wr_en_mem2_16,
  input          io_wr_en_mem2_17,
  input          io_wr_en_mem2_18,
  input          io_wr_en_mem2_19,
  input          io_wr_en_mem2_20,
  input          io_wr_en_mem3_0,
  input          io_wr_en_mem3_1,
  input          io_wr_en_mem3_2,
  input          io_wr_en_mem3_3,
  input          io_wr_en_mem3_4,
  input          io_wr_en_mem3_5,
  input          io_wr_en_mem3_6,
  input          io_wr_en_mem3_7,
  input          io_wr_en_mem3_8,
  input          io_wr_en_mem3_9,
  input          io_wr_en_mem3_10,
  input          io_wr_en_mem3_11,
  input          io_wr_en_mem3_12,
  input          io_wr_en_mem3_13,
  input          io_wr_en_mem3_14,
  input          io_wr_en_mem3_15,
  input          io_wr_en_mem3_16,
  input          io_wr_en_mem3_17,
  input          io_wr_en_mem3_18,
  input          io_wr_en_mem3_19,
  input          io_wr_en_mem3_20,
  input          io_wr_en_mem4_0,
  input          io_wr_en_mem4_1,
  input          io_wr_en_mem4_2,
  input          io_wr_en_mem4_3,
  input          io_wr_en_mem4_4,
  input          io_wr_en_mem4_5,
  input          io_wr_en_mem4_6,
  input          io_wr_en_mem4_7,
  input          io_wr_en_mem4_8,
  input          io_wr_en_mem4_9,
  input          io_wr_en_mem4_10,
  input          io_wr_en_mem4_11,
  input          io_wr_en_mem4_12,
  input          io_wr_en_mem4_13,
  input          io_wr_en_mem4_14,
  input          io_wr_en_mem4_15,
  input          io_wr_en_mem4_16,
  input          io_wr_en_mem4_17,
  input          io_wr_en_mem4_18,
  input          io_wr_en_mem4_19,
  input          io_wr_en_mem4_20,
  input          io_wr_en_mem5_0,
  input          io_wr_en_mem5_1,
  input          io_wr_en_mem5_2,
  input          io_wr_en_mem5_3,
  input          io_wr_en_mem5_4,
  input          io_wr_en_mem5_5,
  input          io_wr_en_mem5_6,
  input          io_wr_en_mem5_7,
  input          io_wr_en_mem5_8,
  input          io_wr_en_mem5_9,
  input          io_wr_en_mem5_10,
  input          io_wr_en_mem5_11,
  input          io_wr_en_mem5_12,
  input          io_wr_en_mem5_13,
  input          io_wr_en_mem5_14,
  input          io_wr_en_mem5_15,
  input          io_wr_en_mem5_16,
  input          io_wr_en_mem5_17,
  input          io_wr_en_mem5_18,
  input          io_wr_en_mem5_19,
  input          io_wr_en_mem5_20,
  input          io_wr_en_mem6_0,
  input          io_wr_en_mem6_1,
  input          io_wr_en_mem6_2,
  input          io_wr_en_mem6_3,
  input          io_wr_en_mem6_4,
  input          io_wr_en_mem6_5,
  input          io_wr_en_mem6_6,
  input          io_wr_en_mem6_7,
  input          io_wr_en_mem6_8,
  input          io_wr_en_mem6_9,
  input          io_wr_en_mem6_10,
  input          io_wr_en_mem6_11,
  input          io_wr_en_mem6_12,
  input          io_wr_en_mem6_13,
  input          io_wr_en_mem6_14,
  input          io_wr_en_mem6_15,
  input          io_wr_en_mem6_16,
  input          io_wr_en_mem6_17,
  input          io_wr_en_mem6_18,
  input          io_wr_en_mem6_19,
  input          io_wr_en_mem6_20,
  input  [287:0] io_wr_instr_mem1_0,
  input  [287:0] io_wr_instr_mem1_1,
  input  [287:0] io_wr_instr_mem1_2,
  input  [287:0] io_wr_instr_mem1_3,
  input  [287:0] io_wr_instr_mem1_4,
  input  [287:0] io_wr_instr_mem1_5,
  input  [287:0] io_wr_instr_mem1_6,
  input  [287:0] io_wr_instr_mem1_7,
  input  [287:0] io_wr_instr_mem1_8,
  input  [287:0] io_wr_instr_mem1_9,
  input  [287:0] io_wr_instr_mem1_10,
  input  [287:0] io_wr_instr_mem1_11,
  input  [287:0] io_wr_instr_mem1_12,
  input  [287:0] io_wr_instr_mem1_13,
  input  [287:0] io_wr_instr_mem1_14,
  input  [287:0] io_wr_instr_mem1_15,
  input  [287:0] io_wr_instr_mem1_16,
  input  [287:0] io_wr_instr_mem1_17,
  input  [287:0] io_wr_instr_mem1_18,
  input  [287:0] io_wr_instr_mem1_19,
  input  [287:0] io_wr_instr_mem1_20,
  input  [127:0] io_wr_instr_mem2_0,
  input  [127:0] io_wr_instr_mem2_1,
  input  [127:0] io_wr_instr_mem2_2,
  input  [127:0] io_wr_instr_mem2_3,
  input  [127:0] io_wr_instr_mem2_4,
  input  [127:0] io_wr_instr_mem2_5,
  input  [127:0] io_wr_instr_mem2_6,
  input  [127:0] io_wr_instr_mem2_7,
  input  [127:0] io_wr_instr_mem2_8,
  input  [127:0] io_wr_instr_mem2_9,
  input  [127:0] io_wr_instr_mem2_10,
  input  [127:0] io_wr_instr_mem2_11,
  input  [127:0] io_wr_instr_mem2_12,
  input  [127:0] io_wr_instr_mem2_13,
  input  [127:0] io_wr_instr_mem2_14,
  input  [127:0] io_wr_instr_mem2_15,
  input  [127:0] io_wr_instr_mem2_16,
  input  [127:0] io_wr_instr_mem2_17,
  input  [127:0] io_wr_instr_mem2_18,
  input  [127:0] io_wr_instr_mem2_19,
  input  [127:0] io_wr_instr_mem2_20,
  input  [127:0] io_wr_instr_mem3_0,
  input  [127:0] io_wr_instr_mem3_1,
  input  [127:0] io_wr_instr_mem3_2,
  input  [127:0] io_wr_instr_mem3_3,
  input  [127:0] io_wr_instr_mem3_4,
  input  [127:0] io_wr_instr_mem3_5,
  input  [127:0] io_wr_instr_mem3_6,
  input  [127:0] io_wr_instr_mem3_7,
  input  [127:0] io_wr_instr_mem3_8,
  input  [127:0] io_wr_instr_mem3_9,
  input  [127:0] io_wr_instr_mem3_10,
  input  [127:0] io_wr_instr_mem3_11,
  input  [127:0] io_wr_instr_mem3_12,
  input  [127:0] io_wr_instr_mem3_13,
  input  [127:0] io_wr_instr_mem3_14,
  input  [127:0] io_wr_instr_mem3_15,
  input  [127:0] io_wr_instr_mem3_16,
  input  [127:0] io_wr_instr_mem3_17,
  input  [127:0] io_wr_instr_mem3_18,
  input  [127:0] io_wr_instr_mem3_19,
  input  [127:0] io_wr_instr_mem3_20,
  input  [127:0] io_wr_instr_mem4_0,
  input  [127:0] io_wr_instr_mem4_1,
  input  [127:0] io_wr_instr_mem4_2,
  input  [127:0] io_wr_instr_mem4_3,
  input  [127:0] io_wr_instr_mem4_4,
  input  [127:0] io_wr_instr_mem4_5,
  input  [127:0] io_wr_instr_mem4_6,
  input  [127:0] io_wr_instr_mem4_7,
  input  [127:0] io_wr_instr_mem4_8,
  input  [127:0] io_wr_instr_mem4_9,
  input  [127:0] io_wr_instr_mem4_10,
  input  [127:0] io_wr_instr_mem4_11,
  input  [127:0] io_wr_instr_mem4_12,
  input  [127:0] io_wr_instr_mem4_13,
  input  [127:0] io_wr_instr_mem4_14,
  input  [127:0] io_wr_instr_mem4_15,
  input  [127:0] io_wr_instr_mem4_16,
  input  [127:0] io_wr_instr_mem4_17,
  input  [127:0] io_wr_instr_mem4_18,
  input  [127:0] io_wr_instr_mem4_19,
  input  [127:0] io_wr_instr_mem4_20,
  input  [127:0] io_wr_instr_mem5_0,
  input  [127:0] io_wr_instr_mem5_1,
  input  [127:0] io_wr_instr_mem5_2,
  input  [127:0] io_wr_instr_mem5_3,
  input  [127:0] io_wr_instr_mem5_4,
  input  [127:0] io_wr_instr_mem5_5,
  input  [127:0] io_wr_instr_mem5_6,
  input  [127:0] io_wr_instr_mem5_7,
  input  [127:0] io_wr_instr_mem5_8,
  input  [127:0] io_wr_instr_mem5_9,
  input  [127:0] io_wr_instr_mem5_10,
  input  [127:0] io_wr_instr_mem5_11,
  input  [127:0] io_wr_instr_mem5_12,
  input  [127:0] io_wr_instr_mem5_13,
  input  [127:0] io_wr_instr_mem5_14,
  input  [127:0] io_wr_instr_mem5_15,
  input  [127:0] io_wr_instr_mem5_16,
  input  [127:0] io_wr_instr_mem5_17,
  input  [127:0] io_wr_instr_mem5_18,
  input  [127:0] io_wr_instr_mem5_19,
  input  [127:0] io_wr_instr_mem5_20,
  input  [127:0] io_wr_instr_mem6_0,
  input  [127:0] io_wr_instr_mem6_1,
  input  [127:0] io_wr_instr_mem6_2,
  input  [127:0] io_wr_instr_mem6_3,
  input  [127:0] io_wr_instr_mem6_4,
  input  [127:0] io_wr_instr_mem6_5,
  input  [127:0] io_wr_instr_mem6_6,
  input  [127:0] io_wr_instr_mem6_7,
  input  [127:0] io_wr_instr_mem6_8,
  input  [127:0] io_wr_instr_mem6_9,
  input  [127:0] io_wr_instr_mem6_10,
  input  [127:0] io_wr_instr_mem6_11,
  input  [127:0] io_wr_instr_mem6_12,
  input  [127:0] io_wr_instr_mem6_13,
  input  [127:0] io_wr_instr_mem6_14,
  input  [127:0] io_wr_instr_mem6_15,
  input  [127:0] io_wr_instr_mem6_16,
  input  [127:0] io_wr_instr_mem6_17,
  input  [127:0] io_wr_instr_mem6_18,
  input  [127:0] io_wr_instr_mem6_19,
  input  [127:0] io_wr_instr_mem6_20,
  input          io_beginRun,
  input          io_wr_D_inBuf_0_validBit,
  input  [3:0]   io_wr_D_inBuf_0_data,
  input          io_wr_D_inBuf_1_validBit,
  input  [3:0]   io_wr_D_inBuf_1_data,
  input          io_wr_D_inBuf_2_validBit,
  input  [3:0]   io_wr_D_inBuf_2_data,
  input          io_wr_D_inBuf_3_validBit,
  input  [3:0]   io_wr_D_inBuf_3_data,
  input          io_wr_D_inBuf_4_validBit,
  input  [3:0]   io_wr_D_inBuf_4_data,
  input          io_wr_D_inBuf_5_validBit,
  input  [3:0]   io_wr_D_inBuf_5_data,
  input          io_wr_D_inBuf_6_validBit,
  input  [3:0]   io_wr_D_inBuf_6_data,
  input          io_wr_D_inBuf_7_validBit,
  input  [3:0]   io_wr_D_inBuf_7_data,
  input          io_wr_D_inBuf_8_validBit,
  input  [3:0]   io_wr_D_inBuf_8_data,
  input          io_wr_D_inBuf_9_validBit,
  input  [3:0]   io_wr_D_inBuf_9_data,
  input          io_wr_D_inBuf_10_validBit,
  input  [3:0]   io_wr_D_inBuf_10_data,
  input          io_wr_D_inBuf_11_validBit,
  input  [3:0]   io_wr_D_inBuf_11_data,
  input          io_wr_D_inBuf_12_validBit,
  input  [3:0]   io_wr_D_inBuf_12_data,
  input          io_wr_D_inBuf_13_validBit,
  input  [3:0]   io_wr_D_inBuf_13_data,
  input          io_wr_D_inBuf_14_validBit,
  input  [3:0]   io_wr_D_inBuf_14_data,
  input          io_wr_D_inBuf_15_validBit,
  input  [3:0]   io_wr_D_inBuf_15_data,
  input          io_wr_D_inBuf_16_validBit,
  input  [3:0]   io_wr_D_inBuf_16_data,
  input          io_wr_D_inBuf_17_validBit,
  input  [3:0]   io_wr_D_inBuf_17_data,
  input          io_wr_D_inBuf_18_validBit,
  input  [3:0]   io_wr_D_inBuf_18_data,
  input          io_wr_D_inBuf_19_validBit,
  input  [3:0]   io_wr_D_inBuf_19_data,
  input          io_wr_D_inBuf_20_validBit,
  input  [3:0]   io_wr_D_inBuf_20_data,
  input          io_wr_D_inBuf_21_validBit,
  input  [3:0]   io_wr_D_inBuf_21_data,
  input          io_wr_D_inBuf_22_validBit,
  input  [3:0]   io_wr_D_inBuf_22_data,
  input          io_wr_D_inBuf_23_validBit,
  input  [3:0]   io_wr_D_inBuf_23_data,
  input          io_wr_D_inBuf_24_validBit,
  input  [3:0]   io_wr_D_inBuf_24_data,
  input          io_wr_D_inBuf_25_validBit,
  input  [3:0]   io_wr_D_inBuf_25_data,
  input          io_wr_D_inBuf_26_validBit,
  input  [3:0]   io_wr_D_inBuf_26_data,
  input          io_wr_D_inBuf_27_validBit,
  input  [3:0]   io_wr_D_inBuf_27_data,
  input          io_wr_D_inBuf_28_validBit,
  input  [3:0]   io_wr_D_inBuf_28_data,
  input          io_wr_D_inBuf_29_validBit,
  input  [3:0]   io_wr_D_inBuf_29_data,
  input          io_wr_D_inBuf_30_validBit,
  input  [3:0]   io_wr_D_inBuf_30_data,
  input          io_wr_D_inBuf_31_validBit,
  input  [3:0]   io_wr_D_inBuf_31_data,
  input          io_wr_D_inBuf_32_validBit,
  input  [3:0]   io_wr_D_inBuf_32_data,
  input          io_wr_D_inBuf_33_validBit,
  input  [3:0]   io_wr_D_inBuf_33_data,
  input          io_wr_D_inBuf_34_validBit,
  input  [3:0]   io_wr_D_inBuf_34_data,
  input          io_wr_D_inBuf_35_validBit,
  input  [3:0]   io_wr_D_inBuf_35_data,
  input          io_wr_D_inBuf_36_validBit,
  input  [3:0]   io_wr_D_inBuf_36_data,
  input          io_wr_D_inBuf_37_validBit,
  input  [3:0]   io_wr_D_inBuf_37_data,
  input          io_wr_D_inBuf_38_validBit,
  input  [3:0]   io_wr_D_inBuf_38_data,
  input          io_wr_D_inBuf_39_validBit,
  input  [3:0]   io_wr_D_inBuf_39_data,
  input          io_wr_D_inBuf_40_validBit,
  input  [3:0]   io_wr_D_inBuf_40_data,
  input          io_wr_D_inBuf_41_validBit,
  input  [3:0]   io_wr_D_inBuf_41_data,
  input          io_wr_D_inBuf_42_validBit,
  input  [3:0]   io_wr_D_inBuf_42_data,
  input          io_wr_D_inBuf_43_validBit,
  input  [3:0]   io_wr_D_inBuf_43_data,
  input          io_wr_D_inBuf_44_validBit,
  input  [3:0]   io_wr_D_inBuf_44_data,
  input          io_wr_D_inBuf_45_validBit,
  input  [3:0]   io_wr_D_inBuf_45_data,
  input          io_wr_D_inBuf_46_validBit,
  input  [3:0]   io_wr_D_inBuf_46_data,
  input          io_wr_D_inBuf_47_validBit,
  input  [3:0]   io_wr_D_inBuf_47_data,
  input          io_wr_D_inBuf_48_validBit,
  input  [3:0]   io_wr_D_inBuf_48_data,
  input          io_wr_D_inBuf_49_validBit,
  input  [3:0]   io_wr_D_inBuf_49_data,
  input          io_wr_D_inBuf_50_validBit,
  input  [3:0]   io_wr_D_inBuf_50_data,
  input          io_wr_D_inBuf_51_validBit,
  input  [3:0]   io_wr_D_inBuf_51_data,
  input          io_wr_D_inBuf_52_validBit,
  input  [3:0]   io_wr_D_inBuf_52_data,
  input          io_wr_D_inBuf_53_validBit,
  input  [3:0]   io_wr_D_inBuf_53_data,
  input          io_wr_D_inBuf_54_validBit,
  input  [3:0]   io_wr_D_inBuf_54_data,
  input          io_wr_D_inBuf_55_validBit,
  input  [3:0]   io_wr_D_inBuf_55_data,
  input          io_wr_D_inBuf_56_validBit,
  input  [3:0]   io_wr_D_inBuf_56_data,
  input          io_wr_D_inBuf_57_validBit,
  input  [3:0]   io_wr_D_inBuf_57_data,
  input          io_wr_D_inBuf_58_validBit,
  input  [3:0]   io_wr_D_inBuf_58_data,
  input          io_wr_D_inBuf_59_validBit,
  input  [3:0]   io_wr_D_inBuf_59_data,
  input          io_wr_D_inBuf_60_validBit,
  input  [3:0]   io_wr_D_inBuf_60_data,
  input          io_wr_D_inBuf_61_validBit,
  input  [3:0]   io_wr_D_inBuf_61_data,
  input          io_wr_D_inBuf_62_validBit,
  input  [3:0]   io_wr_D_inBuf_62_data,
  input          io_wr_D_inBuf_63_validBit,
  input  [3:0]   io_wr_D_inBuf_63_data,
  input  [1:0]   io_wr_Tag_inBuf,
  input          io_wr_Addr_inBuf_en,
  input  [7:0]   io_rd_Addr_outBuf,
  output         io_rd_D_outBuf_0_validBit,
  output [3:0]   io_rd_D_outBuf_0_data,
  output         io_rd_D_outBuf_1_validBit,
  output [3:0]   io_rd_D_outBuf_1_data,
  output         io_rd_D_outBuf_2_validBit,
  output [3:0]   io_rd_D_outBuf_2_data,
  output         io_rd_D_outBuf_3_validBit,
  output [3:0]   io_rd_D_outBuf_3_data,
  output         io_rd_D_outBuf_4_validBit,
  output [3:0]   io_rd_D_outBuf_4_data,
  output         io_rd_D_outBuf_5_validBit,
  output [3:0]   io_rd_D_outBuf_5_data,
  output         io_rd_D_outBuf_6_validBit,
  output [3:0]   io_rd_D_outBuf_6_data,
  output         io_rd_D_outBuf_7_validBit,
  output [3:0]   io_rd_D_outBuf_7_data,
  output         io_rd_D_outBuf_8_validBit,
  output [3:0]   io_rd_D_outBuf_8_data,
  output         io_rd_D_outBuf_9_validBit,
  output [3:0]   io_rd_D_outBuf_9_data,
  output         io_rd_D_outBuf_10_validBit,
  output [3:0]   io_rd_D_outBuf_10_data,
  output         io_rd_D_outBuf_11_validBit,
  output [3:0]   io_rd_D_outBuf_11_data,
  output         io_rd_D_outBuf_12_validBit,
  output [3:0]   io_rd_D_outBuf_12_data,
  output         io_rd_D_outBuf_13_validBit,
  output [3:0]   io_rd_D_outBuf_13_data,
  output         io_rd_D_outBuf_14_validBit,
  output [3:0]   io_rd_D_outBuf_14_data,
  output         io_rd_D_outBuf_15_validBit,
  output [3:0]   io_rd_D_outBuf_15_data,
  output         io_rd_D_outBuf_16_validBit,
  output [3:0]   io_rd_D_outBuf_16_data,
  output         io_rd_D_outBuf_17_validBit,
  output [3:0]   io_rd_D_outBuf_17_data,
  output         io_rd_D_outBuf_18_validBit,
  output [3:0]   io_rd_D_outBuf_18_data,
  output         io_rd_D_outBuf_19_validBit,
  output [3:0]   io_rd_D_outBuf_19_data,
  output         io_rd_D_outBuf_20_validBit,
  output [3:0]   io_rd_D_outBuf_20_data,
  output         io_rd_D_outBuf_21_validBit,
  output [3:0]   io_rd_D_outBuf_21_data,
  output         io_rd_D_outBuf_22_validBit,
  output [3:0]   io_rd_D_outBuf_22_data,
  output         io_rd_D_outBuf_23_validBit,
  output [3:0]   io_rd_D_outBuf_23_data,
  output         io_rd_D_outBuf_24_validBit,
  output [3:0]   io_rd_D_outBuf_24_data,
  output         io_rd_D_outBuf_25_validBit,
  output [3:0]   io_rd_D_outBuf_25_data,
  output         io_rd_D_outBuf_26_validBit,
  output [3:0]   io_rd_D_outBuf_26_data,
  output         io_rd_D_outBuf_27_validBit,
  output [3:0]   io_rd_D_outBuf_27_data,
  output         io_rd_D_outBuf_28_validBit,
  output [3:0]   io_rd_D_outBuf_28_data,
  output         io_rd_D_outBuf_29_validBit,
  output [3:0]   io_rd_D_outBuf_29_data,
  output         io_rd_D_outBuf_30_validBit,
  output [3:0]   io_rd_D_outBuf_30_data,
  output         io_rd_D_outBuf_31_validBit,
  output [3:0]   io_rd_D_outBuf_31_data,
  output         io_rd_D_outBuf_32_validBit,
  output [3:0]   io_rd_D_outBuf_32_data,
  output         io_rd_D_outBuf_33_validBit,
  output [3:0]   io_rd_D_outBuf_33_data,
  output         io_rd_D_outBuf_34_validBit,
  output [3:0]   io_rd_D_outBuf_34_data,
  output         io_rd_D_outBuf_35_validBit,
  output [3:0]   io_rd_D_outBuf_35_data,
  output         io_rd_D_outBuf_36_validBit,
  output [3:0]   io_rd_D_outBuf_36_data,
  output         io_rd_D_outBuf_37_validBit,
  output [3:0]   io_rd_D_outBuf_37_data,
  output         io_rd_D_outBuf_38_validBit,
  output [3:0]   io_rd_D_outBuf_38_data,
  output         io_rd_D_outBuf_39_validBit,
  output [3:0]   io_rd_D_outBuf_39_data,
  output         io_rd_D_outBuf_40_validBit,
  output [3:0]   io_rd_D_outBuf_40_data,
  output         io_rd_D_outBuf_41_validBit,
  output [3:0]   io_rd_D_outBuf_41_data,
  output         io_rd_D_outBuf_42_validBit,
  output [3:0]   io_rd_D_outBuf_42_data,
  output         io_rd_D_outBuf_43_validBit,
  output [3:0]   io_rd_D_outBuf_43_data,
  output         io_rd_D_outBuf_44_validBit,
  output [3:0]   io_rd_D_outBuf_44_data,
  output         io_rd_D_outBuf_45_validBit,
  output [3:0]   io_rd_D_outBuf_45_data,
  output         io_rd_D_outBuf_46_validBit,
  output [3:0]   io_rd_D_outBuf_46_data,
  output         io_rd_D_outBuf_47_validBit,
  output [3:0]   io_rd_D_outBuf_47_data,
  output         io_rd_D_outBuf_48_validBit,
  output [3:0]   io_rd_D_outBuf_48_data,
  output         io_rd_D_outBuf_49_validBit,
  output [3:0]   io_rd_D_outBuf_49_data,
  output         io_rd_D_outBuf_50_validBit,
  output [3:0]   io_rd_D_outBuf_50_data,
  output         io_rd_D_outBuf_51_validBit,
  output [3:0]   io_rd_D_outBuf_51_data,
  output         io_rd_D_outBuf_52_validBit,
  output [3:0]   io_rd_D_outBuf_52_data,
  output         io_rd_D_outBuf_53_validBit,
  output [3:0]   io_rd_D_outBuf_53_data,
  output         io_rd_D_outBuf_54_validBit,
  output [3:0]   io_rd_D_outBuf_54_data,
  output         io_rd_D_outBuf_55_validBit,
  output [3:0]   io_rd_D_outBuf_55_data,
  output         io_rd_D_outBuf_56_validBit,
  output [3:0]   io_rd_D_outBuf_56_data,
  output         io_rd_D_outBuf_57_validBit,
  output [3:0]   io_rd_D_outBuf_57_data,
  output         io_rd_D_outBuf_58_validBit,
  output [3:0]   io_rd_D_outBuf_58_data,
  output         io_rd_D_outBuf_59_validBit,
  output [3:0]   io_rd_D_outBuf_59_data,
  output         io_rd_D_outBuf_60_validBit,
  output [3:0]   io_rd_D_outBuf_60_data,
  output         io_rd_D_outBuf_61_validBit,
  output [3:0]   io_rd_D_outBuf_61_data,
  output         io_rd_D_outBuf_62_validBit,
  output [3:0]   io_rd_D_outBuf_62_data,
  output         io_rd_D_outBuf_63_validBit,
  output [3:0]   io_rd_D_outBuf_63_data,
  output [7:0]   io_PC_out
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_234;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_261;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_273;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_294;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_300;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_333;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_339;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_345;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_351;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_372;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_378;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_384;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_390;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_398;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_404;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_410;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_416;
  reg [31:0] _RAND_418;
  reg [31:0] _RAND_420;
  reg [31:0] _RAND_422;
  reg [31:0] _RAND_424;
  reg [31:0] _RAND_426;
  reg [31:0] _RAND_428;
  reg [31:0] _RAND_430;
  reg [31:0] _RAND_432;
  reg [31:0] _RAND_434;
  reg [31:0] _RAND_436;
  reg [31:0] _RAND_438;
  reg [31:0] _RAND_440;
  reg [31:0] _RAND_442;
  reg [31:0] _RAND_444;
  reg [31:0] _RAND_446;
  reg [31:0] _RAND_448;
  reg [31:0] _RAND_450;
  reg [31:0] _RAND_452;
  reg [31:0] _RAND_454;
  reg [31:0] _RAND_456;
  reg [31:0] _RAND_458;
  reg [31:0] _RAND_460;
  reg [31:0] _RAND_462;
  reg [31:0] _RAND_464;
  reg [31:0] _RAND_466;
  reg [31:0] _RAND_468;
  reg [31:0] _RAND_470;
  reg [31:0] _RAND_472;
  reg [31:0] _RAND_474;
  reg [31:0] _RAND_476;
  reg [31:0] _RAND_478;
  reg [31:0] _RAND_480;
  reg [31:0] _RAND_482;
  reg [31:0] _RAND_484;
  reg [31:0] _RAND_486;
  reg [31:0] _RAND_488;
  reg [31:0] _RAND_490;
  reg [31:0] _RAND_492;
  reg [31:0] _RAND_494;
  reg [31:0] _RAND_496;
  reg [31:0] _RAND_498;
  reg [31:0] _RAND_500;
  reg [31:0] _RAND_502;
  reg [31:0] _RAND_504;
  reg [31:0] _RAND_506;
  reg [31:0] _RAND_508;
  reg [31:0] _RAND_510;
  reg [31:0] _RAND_512;
  reg [31:0] _RAND_514;
  reg [31:0] _RAND_516;
  reg [31:0] _RAND_518;
  reg [31:0] _RAND_520;
  reg [31:0] _RAND_522;
  reg [31:0] _RAND_524;
  reg [31:0] _RAND_526;
  reg [31:0] _RAND_528;
  reg [31:0] _RAND_530;
  reg [31:0] _RAND_532;
  reg [31:0] _RAND_534;
  reg [31:0] _RAND_536;
  reg [31:0] _RAND_538;
  reg [31:0] _RAND_540;
  reg [31:0] _RAND_542;
  reg [31:0] _RAND_544;
  reg [31:0] _RAND_546;
  reg [31:0] _RAND_548;
  reg [31:0] _RAND_550;
  reg [31:0] _RAND_552;
  reg [31:0] _RAND_554;
  reg [31:0] _RAND_556;
  reg [31:0] _RAND_558;
  reg [31:0] _RAND_560;
  reg [31:0] _RAND_562;
  reg [31:0] _RAND_564;
  reg [31:0] _RAND_566;
  reg [31:0] _RAND_568;
  reg [31:0] _RAND_570;
  reg [31:0] _RAND_572;
  reg [31:0] _RAND_574;
  reg [31:0] _RAND_576;
  reg [31:0] _RAND_578;
  reg [31:0] _RAND_580;
  reg [31:0] _RAND_582;
  reg [31:0] _RAND_584;
  reg [31:0] _RAND_586;
  reg [31:0] _RAND_588;
  reg [31:0] _RAND_590;
  reg [31:0] _RAND_592;
  reg [31:0] _RAND_594;
  reg [31:0] _RAND_596;
  reg [31:0] _RAND_598;
  reg [31:0] _RAND_600;
  reg [31:0] _RAND_602;
  reg [31:0] _RAND_604;
  reg [31:0] _RAND_606;
  reg [31:0] _RAND_608;
  reg [31:0] _RAND_610;
  reg [31:0] _RAND_612;
  reg [31:0] _RAND_614;
  reg [31:0] _RAND_616;
  reg [31:0] _RAND_618;
  reg [31:0] _RAND_620;
  reg [31:0] _RAND_622;
  reg [31:0] _RAND_624;
  reg [31:0] _RAND_626;
  reg [31:0] _RAND_628;
  reg [31:0] _RAND_630;
  reg [31:0] _RAND_632;
  reg [31:0] _RAND_634;
  reg [31:0] _RAND_636;
  reg [31:0] _RAND_638;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_280;
  reg [31:0] _RAND_281;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_319;
  reg [31:0] _RAND_320;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_325;
  reg [31:0] _RAND_326;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_358;
  reg [31:0] _RAND_359;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_364;
  reg [31:0] _RAND_365;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_385;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_391;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_397;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_403;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_411;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_415;
  reg [31:0] _RAND_417;
  reg [31:0] _RAND_419;
  reg [31:0] _RAND_421;
  reg [31:0] _RAND_423;
  reg [31:0] _RAND_425;
  reg [31:0] _RAND_427;
  reg [31:0] _RAND_429;
  reg [31:0] _RAND_431;
  reg [31:0] _RAND_433;
  reg [31:0] _RAND_435;
  reg [31:0] _RAND_437;
  reg [31:0] _RAND_439;
  reg [31:0] _RAND_441;
  reg [31:0] _RAND_443;
  reg [31:0] _RAND_445;
  reg [31:0] _RAND_447;
  reg [31:0] _RAND_449;
  reg [31:0] _RAND_451;
  reg [31:0] _RAND_453;
  reg [31:0] _RAND_455;
  reg [31:0] _RAND_457;
  reg [31:0] _RAND_459;
  reg [31:0] _RAND_461;
  reg [31:0] _RAND_463;
  reg [31:0] _RAND_465;
  reg [31:0] _RAND_467;
  reg [31:0] _RAND_469;
  reg [31:0] _RAND_471;
  reg [31:0] _RAND_473;
  reg [31:0] _RAND_475;
  reg [31:0] _RAND_477;
  reg [31:0] _RAND_479;
  reg [31:0] _RAND_481;
  reg [31:0] _RAND_483;
  reg [31:0] _RAND_485;
  reg [31:0] _RAND_487;
  reg [31:0] _RAND_489;
  reg [31:0] _RAND_491;
  reg [31:0] _RAND_493;
  reg [31:0] _RAND_495;
  reg [31:0] _RAND_497;
  reg [31:0] _RAND_499;
  reg [31:0] _RAND_501;
  reg [31:0] _RAND_503;
  reg [31:0] _RAND_505;
  reg [31:0] _RAND_507;
  reg [31:0] _RAND_509;
  reg [31:0] _RAND_511;
  reg [31:0] _RAND_513;
  reg [31:0] _RAND_515;
  reg [31:0] _RAND_517;
  reg [31:0] _RAND_519;
  reg [31:0] _RAND_521;
  reg [31:0] _RAND_523;
  reg [31:0] _RAND_525;
  reg [31:0] _RAND_527;
  reg [31:0] _RAND_529;
  reg [31:0] _RAND_531;
  reg [31:0] _RAND_533;
  reg [31:0] _RAND_535;
  reg [31:0] _RAND_537;
  reg [31:0] _RAND_539;
  reg [31:0] _RAND_541;
  reg [31:0] _RAND_543;
  reg [31:0] _RAND_545;
  reg [31:0] _RAND_547;
  reg [31:0] _RAND_549;
  reg [31:0] _RAND_551;
  reg [31:0] _RAND_553;
  reg [31:0] _RAND_555;
  reg [31:0] _RAND_557;
  reg [31:0] _RAND_559;
  reg [31:0] _RAND_561;
  reg [31:0] _RAND_563;
  reg [31:0] _RAND_565;
  reg [31:0] _RAND_567;
  reg [31:0] _RAND_569;
  reg [31:0] _RAND_571;
  reg [31:0] _RAND_573;
  reg [31:0] _RAND_575;
  reg [31:0] _RAND_577;
  reg [31:0] _RAND_579;
  reg [31:0] _RAND_581;
  reg [31:0] _RAND_583;
  reg [31:0] _RAND_585;
  reg [31:0] _RAND_587;
  reg [31:0] _RAND_589;
  reg [31:0] _RAND_591;
  reg [31:0] _RAND_593;
  reg [31:0] _RAND_595;
  reg [31:0] _RAND_597;
  reg [31:0] _RAND_599;
  reg [31:0] _RAND_601;
  reg [31:0] _RAND_603;
  reg [31:0] _RAND_605;
  reg [31:0] _RAND_607;
  reg [31:0] _RAND_609;
  reg [31:0] _RAND_611;
  reg [31:0] _RAND_613;
  reg [31:0] _RAND_615;
  reg [31:0] _RAND_617;
  reg [31:0] _RAND_619;
  reg [31:0] _RAND_621;
  reg [31:0] _RAND_623;
  reg [31:0] _RAND_625;
  reg [31:0] _RAND_627;
  reg [31:0] _RAND_629;
  reg [31:0] _RAND_631;
  reg [31:0] _RAND_633;
  reg [31:0] _RAND_635;
  reg [31:0] _RAND_637;
  reg [31:0] _RAND_639;
  reg [31:0] _RAND_640;
  reg [31:0] _RAND_641;
  reg [31:0] _RAND_642;
  reg [31:0] _RAND_643;
  reg [31:0] _RAND_644;
  reg [31:0] _RAND_645;
  reg [31:0] _RAND_646;
  reg [31:0] _RAND_647;
  reg [31:0] _RAND_648;
  reg [31:0] _RAND_649;
  reg [31:0] _RAND_650;
  reg [31:0] _RAND_651;
  reg [31:0] _RAND_652;
  reg [31:0] _RAND_653;
  reg [31:0] _RAND_654;
  reg [31:0] _RAND_655;
  reg [31:0] _RAND_656;
  reg [31:0] _RAND_657;
  reg [31:0] _RAND_658;
  reg [31:0] _RAND_659;
  reg [31:0] _RAND_660;
  reg [31:0] _RAND_661;
  reg [31:0] _RAND_662;
  reg [31:0] _RAND_663;
  reg [31:0] _RAND_664;
  reg [31:0] _RAND_665;
  reg [31:0] _RAND_666;
  reg [31:0] _RAND_667;
  reg [31:0] _RAND_668;
  reg [31:0] _RAND_669;
  reg [31:0] _RAND_670;
  reg [31:0] _RAND_671;
  reg [31:0] _RAND_672;
  reg [31:0] _RAND_673;
  reg [31:0] _RAND_674;
  reg [31:0] _RAND_675;
  reg [31:0] _RAND_676;
  reg [31:0] _RAND_677;
  reg [31:0] _RAND_678;
  reg [31:0] _RAND_679;
  reg [31:0] _RAND_680;
  reg [31:0] _RAND_681;
  reg [31:0] _RAND_682;
  reg [31:0] _RAND_683;
  reg [31:0] _RAND_684;
  reg [31:0] _RAND_685;
  reg [31:0] _RAND_686;
  reg [31:0] _RAND_687;
  reg [31:0] _RAND_688;
  reg [31:0] _RAND_689;
  reg [31:0] _RAND_690;
  reg [31:0] _RAND_691;
  reg [31:0] _RAND_692;
  reg [31:0] _RAND_693;
  reg [31:0] _RAND_694;
  reg [31:0] _RAND_695;
  reg [31:0] _RAND_696;
  reg [31:0] _RAND_697;
  reg [31:0] _RAND_698;
  reg [31:0] _RAND_699;
  reg [31:0] _RAND_700;
  reg [31:0] _RAND_701;
  reg [31:0] _RAND_702;
  reg [31:0] _RAND_703;
  reg [31:0] _RAND_704;
  reg [31:0] _RAND_705;
  reg [31:0] _RAND_706;
  reg [31:0] _RAND_707;
  reg [31:0] _RAND_708;
  reg [31:0] _RAND_709;
  reg [31:0] _RAND_710;
  reg [31:0] _RAND_711;
  reg [31:0] _RAND_712;
  reg [31:0] _RAND_713;
  reg [31:0] _RAND_714;
  reg [31:0] _RAND_715;
  reg [31:0] _RAND_716;
  reg [31:0] _RAND_717;
  reg [31:0] _RAND_718;
  reg [31:0] _RAND_719;
  reg [31:0] _RAND_720;
  reg [31:0] _RAND_721;
  reg [31:0] _RAND_722;
  reg [31:0] _RAND_723;
  reg [31:0] _RAND_724;
  reg [31:0] _RAND_725;
  reg [31:0] _RAND_726;
  reg [31:0] _RAND_727;
  reg [31:0] _RAND_728;
  reg [31:0] _RAND_729;
  reg [31:0] _RAND_730;
  reg [31:0] _RAND_731;
  reg [31:0] _RAND_732;
  reg [31:0] _RAND_733;
  reg [31:0] _RAND_734;
  reg [31:0] _RAND_735;
  reg [31:0] _RAND_736;
  reg [31:0] _RAND_737;
  reg [31:0] _RAND_738;
  reg [31:0] _RAND_739;
  reg [31:0] _RAND_740;
  reg [31:0] _RAND_741;
  reg [31:0] _RAND_742;
  reg [31:0] _RAND_743;
  reg [31:0] _RAND_744;
  reg [31:0] _RAND_745;
  reg [31:0] _RAND_746;
  reg [31:0] _RAND_747;
  reg [31:0] _RAND_748;
  reg [31:0] _RAND_749;
  reg [31:0] _RAND_750;
  reg [31:0] _RAND_751;
  reg [31:0] _RAND_752;
  reg [31:0] _RAND_753;
  reg [31:0] _RAND_754;
  reg [31:0] _RAND_755;
  reg [31:0] _RAND_756;
  reg [31:0] _RAND_757;
  reg [31:0] _RAND_758;
  reg [31:0] _RAND_759;
  reg [31:0] _RAND_760;
  reg [31:0] _RAND_761;
  reg [31:0] _RAND_762;
  reg [31:0] _RAND_763;
  reg [31:0] _RAND_764;
  reg [31:0] _RAND_765;
  reg [31:0] _RAND_766;
  reg [31:0] _RAND_767;
  reg [31:0] _RAND_768;
  reg [31:0] _RAND_769;
  reg [31:0] _RAND_770;
  reg [31:0] _RAND_771;
  reg [31:0] _RAND_772;
  reg [31:0] _RAND_773;
  reg [31:0] _RAND_774;
  reg [31:0] _RAND_775;
  reg [31:0] _RAND_776;
  reg [31:0] _RAND_777;
  reg [31:0] _RAND_778;
  reg [31:0] _RAND_779;
  reg [31:0] _RAND_780;
  reg [31:0] _RAND_781;
  reg [31:0] _RAND_782;
  reg [31:0] _RAND_783;
  reg [31:0] _RAND_784;
  reg [31:0] _RAND_785;
  reg [31:0] _RAND_786;
  reg [31:0] _RAND_787;
  reg [31:0] _RAND_788;
  reg [31:0] _RAND_789;
  reg [31:0] _RAND_790;
  reg [31:0] _RAND_791;
  reg [31:0] _RAND_792;
  reg [31:0] _RAND_793;
  reg [31:0] _RAND_794;
  reg [31:0] _RAND_795;
  reg [31:0] _RAND_796;
  reg [31:0] _RAND_797;
  reg [31:0] _RAND_798;
  reg [31:0] _RAND_799;
  reg [31:0] _RAND_800;
  reg [31:0] _RAND_801;
  reg [31:0] _RAND_802;
  reg [31:0] _RAND_803;
  reg [31:0] _RAND_804;
  reg [31:0] _RAND_805;
  reg [31:0] _RAND_806;
  reg [31:0] _RAND_807;
  reg [31:0] _RAND_808;
  reg [31:0] _RAND_809;
  reg [31:0] _RAND_810;
  reg [31:0] _RAND_811;
  reg [31:0] _RAND_812;
  reg [31:0] _RAND_813;
  reg [31:0] _RAND_814;
  reg [31:0] _RAND_815;
  reg [31:0] _RAND_816;
  reg [31:0] _RAND_817;
  reg [31:0] _RAND_818;
  reg [31:0] _RAND_819;
  reg [31:0] _RAND_820;
  reg [31:0] _RAND_821;
  reg [31:0] _RAND_822;
  reg [31:0] _RAND_823;
  reg [31:0] _RAND_824;
  reg [31:0] _RAND_825;
  reg [31:0] _RAND_826;
  reg [31:0] _RAND_827;
  reg [31:0] _RAND_828;
  reg [31:0] _RAND_829;
  reg [31:0] _RAND_830;
  reg [31:0] _RAND_831;
  reg [31:0] _RAND_832;
  reg [31:0] _RAND_833;
  reg [31:0] _RAND_834;
  reg [31:0] _RAND_835;
  reg [31:0] _RAND_836;
  reg [31:0] _RAND_837;
  reg [31:0] _RAND_838;
  reg [31:0] _RAND_839;
  reg [31:0] _RAND_840;
  reg [31:0] _RAND_841;
  reg [31:0] _RAND_842;
  reg [31:0] _RAND_843;
  reg [31:0] _RAND_844;
  reg [31:0] _RAND_845;
  reg [31:0] _RAND_846;
  reg [31:0] _RAND_847;
  reg [31:0] _RAND_848;
  reg [31:0] _RAND_849;
  reg [31:0] _RAND_850;
  reg [31:0] _RAND_851;
  reg [31:0] _RAND_852;
  reg [31:0] _RAND_853;
  reg [31:0] _RAND_854;
  reg [31:0] _RAND_855;
  reg [31:0] _RAND_856;
  reg [31:0] _RAND_857;
  reg [31:0] _RAND_858;
  reg [31:0] _RAND_859;
  reg [31:0] _RAND_860;
  reg [31:0] _RAND_861;
  reg [31:0] _RAND_862;
  reg [31:0] _RAND_863;
  reg [31:0] _RAND_864;
  reg [31:0] _RAND_865;
  reg [31:0] _RAND_866;
  reg [31:0] _RAND_867;
  reg [31:0] _RAND_868;
  reg [31:0] _RAND_869;
  reg [31:0] _RAND_870;
  reg [31:0] _RAND_871;
  reg [31:0] _RAND_872;
  reg [31:0] _RAND_873;
  reg [31:0] _RAND_874;
  reg [31:0] _RAND_875;
  reg [31:0] _RAND_876;
  reg [31:0] _RAND_877;
  reg [31:0] _RAND_878;
  reg [31:0] _RAND_879;
  reg [31:0] _RAND_880;
  reg [31:0] _RAND_881;
  reg [31:0] _RAND_882;
  reg [31:0] _RAND_883;
  reg [31:0] _RAND_884;
  reg [31:0] _RAND_885;
  reg [31:0] _RAND_886;
  reg [31:0] _RAND_887;
  reg [31:0] _RAND_888;
  reg [31:0] _RAND_889;
  reg [31:0] _RAND_890;
  reg [31:0] _RAND_891;
  reg [31:0] _RAND_892;
  reg [31:0] _RAND_893;
  reg [31:0] _RAND_894;
  reg [31:0] _RAND_895;
  reg [31:0] _RAND_896;
  reg [31:0] _RAND_897;
  reg [31:0] _RAND_898;
  reg [31:0] _RAND_899;
  reg [31:0] _RAND_900;
`endif // RANDOMIZE_REG_INIT
  reg  inputDataBuffer_0_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_0_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_0_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_0_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_0_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_0_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_0_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_0_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_0_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_0_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_0_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_0_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_0_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_0_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_0_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_0_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_0_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_0_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_1_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_1_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_1_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_1_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_1_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_1_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_1_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_1_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_1_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_1_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_1_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_1_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_1_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_1_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_1_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_1_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_1_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_1_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_2_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_2_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_2_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_2_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_2_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_2_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_2_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_2_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_2_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_2_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_2_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_2_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_2_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_2_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_2_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_2_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_2_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_2_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_3_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_3_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_3_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_3_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_3_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_3_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_3_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_3_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_3_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_3_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_3_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_3_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_3_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_3_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_3_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_3_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_3_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_3_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_4_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_4_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_4_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_4_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_4_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_4_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_4_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_4_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_4_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_4_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_4_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_4_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_4_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_4_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_4_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_4_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_4_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_4_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_5_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_5_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_5_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_5_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_5_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_5_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_5_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_5_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_5_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_5_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_5_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_5_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_5_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_5_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_5_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_5_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_5_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_5_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_6_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_6_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_6_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_6_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_6_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_6_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_6_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_6_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_6_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_6_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_6_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_6_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_6_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_6_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_6_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_6_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_6_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_6_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_7_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_7_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_7_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_7_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_7_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_7_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_7_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_7_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_7_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_7_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_7_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_7_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_7_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_7_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_7_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_7_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_7_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_7_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_8_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_8_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_8_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_8_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_8_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_8_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_8_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_8_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_8_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_8_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_8_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_8_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_8_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_8_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_8_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_8_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_8_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_8_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_9_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_9_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_9_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_9_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_9_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_9_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_9_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_9_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_9_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_9_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_9_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_9_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_9_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_9_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_9_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_9_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_9_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_9_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_10_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_10_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_10_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_10_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_10_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_10_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_10_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_10_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_10_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_10_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_10_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_10_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_10_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_10_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_10_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_10_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_10_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_10_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_11_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_11_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_11_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_11_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_11_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_11_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_11_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_11_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_11_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_11_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_11_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_11_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_11_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_11_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_11_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_11_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_11_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_11_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_12_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_12_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_12_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_12_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_12_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_12_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_12_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_12_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_12_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_12_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_12_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_12_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_12_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_12_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_12_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_12_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_12_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_12_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_13_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_13_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_13_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_13_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_13_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_13_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_13_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_13_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_13_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_13_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_13_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_13_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_13_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_13_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_13_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_13_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_13_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_13_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_14_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_14_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_14_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_14_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_14_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_14_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_14_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_14_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_14_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_14_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_14_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_14_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_14_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_14_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_14_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_14_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_14_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_14_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_15_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_15_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_15_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_15_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_15_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_15_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_15_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_15_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_15_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_15_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_15_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_15_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_15_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_15_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_15_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_15_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_15_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_15_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_16_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_16_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_16_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_16_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_16_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_16_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_16_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_16_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_16_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_16_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_16_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_16_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_16_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_16_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_16_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_16_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_16_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_16_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_17_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_17_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_17_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_17_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_17_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_17_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_17_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_17_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_17_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_17_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_17_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_17_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_17_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_17_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_17_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_17_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_17_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_17_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_18_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_18_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_18_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_18_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_18_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_18_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_18_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_18_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_18_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_18_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_18_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_18_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_18_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_18_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_18_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_18_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_18_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_18_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_19_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_19_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_19_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_19_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_19_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_19_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_19_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_19_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_19_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_19_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_19_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_19_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_19_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_19_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_19_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_19_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_19_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_19_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_20_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_20_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_20_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_20_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_20_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_20_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_20_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_20_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_20_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_20_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_20_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_20_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_20_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_20_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_20_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_20_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_20_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_20_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_21_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_21_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_21_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_21_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_21_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_21_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_21_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_21_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_21_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_21_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_21_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_21_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_21_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_21_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_21_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_21_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_21_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_21_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_22_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_22_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_22_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_22_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_22_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_22_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_22_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_22_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_22_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_22_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_22_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_22_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_22_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_22_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_22_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_22_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_22_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_22_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_23_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_23_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_23_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_23_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_23_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_23_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_23_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_23_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_23_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_23_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_23_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_23_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_23_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_23_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_23_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_23_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_23_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_23_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_24_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_24_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_24_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_24_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_24_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_24_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_24_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_24_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_24_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_24_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_24_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_24_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_24_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_24_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_24_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_24_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_24_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_24_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_25_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_25_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_25_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_25_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_25_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_25_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_25_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_25_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_25_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_25_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_25_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_25_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_25_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_25_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_25_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_25_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_25_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_25_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_26_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_26_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_26_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_26_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_26_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_26_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_26_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_26_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_26_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_26_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_26_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_26_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_26_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_26_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_26_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_26_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_26_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_26_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_27_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_27_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_27_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_27_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_27_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_27_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_27_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_27_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_27_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_27_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_27_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_27_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_27_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_27_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_27_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_27_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_27_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_27_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_28_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_28_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_28_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_28_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_28_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_28_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_28_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_28_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_28_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_28_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_28_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_28_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_28_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_28_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_28_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_28_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_28_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_28_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_29_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_29_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_29_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_29_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_29_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_29_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_29_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_29_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_29_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_29_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_29_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_29_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_29_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_29_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_29_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_29_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_29_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_29_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_30_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_30_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_30_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_30_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_30_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_30_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_30_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_30_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_30_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_30_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_30_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_30_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_30_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_30_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_30_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_30_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_30_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_30_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_31_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_31_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_31_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_31_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_31_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_31_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_31_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_31_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_31_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_31_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_31_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_31_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_31_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_31_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_31_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_31_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_31_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_31_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_32_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_32_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_32_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_32_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_32_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_32_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_32_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_32_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_32_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_32_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_32_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_32_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_32_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_32_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_32_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_32_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_32_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_32_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_33_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_33_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_33_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_33_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_33_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_33_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_33_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_33_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_33_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_33_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_33_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_33_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_33_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_33_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_33_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_33_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_33_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_33_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_34_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_34_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_34_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_34_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_34_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_34_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_34_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_34_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_34_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_34_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_34_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_34_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_34_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_34_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_34_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_34_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_34_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_34_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_35_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_35_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_35_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_35_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_35_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_35_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_35_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_35_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_35_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_35_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_35_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_35_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_35_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_35_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_35_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_35_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_35_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_35_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_36_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_36_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_36_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_36_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_36_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_36_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_36_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_36_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_36_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_36_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_36_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_36_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_36_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_36_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_36_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_36_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_36_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_36_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_37_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_37_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_37_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_37_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_37_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_37_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_37_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_37_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_37_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_37_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_37_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_37_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_37_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_37_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_37_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_37_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_37_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_37_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_38_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_38_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_38_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_38_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_38_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_38_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_38_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_38_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_38_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_38_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_38_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_38_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_38_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_38_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_38_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_38_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_38_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_38_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_39_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_39_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_39_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_39_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_39_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_39_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_39_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_39_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_39_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_39_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_39_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_39_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_39_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_39_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_39_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_39_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_39_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_39_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_40_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_40_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_40_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_40_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_40_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_40_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_40_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_40_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_40_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_40_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_40_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_40_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_40_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_40_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_40_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_40_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_40_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_40_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_41_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_41_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_41_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_41_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_41_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_41_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_41_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_41_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_41_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_41_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_41_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_41_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_41_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_41_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_41_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_41_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_41_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_41_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_42_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_42_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_42_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_42_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_42_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_42_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_42_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_42_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_42_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_42_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_42_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_42_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_42_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_42_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_42_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_42_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_42_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_42_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_43_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_43_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_43_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_43_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_43_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_43_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_43_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_43_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_43_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_43_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_43_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_43_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_43_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_43_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_43_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_43_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_43_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_43_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_44_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_44_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_44_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_44_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_44_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_44_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_44_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_44_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_44_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_44_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_44_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_44_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_44_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_44_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_44_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_44_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_44_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_44_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_45_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_45_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_45_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_45_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_45_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_45_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_45_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_45_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_45_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_45_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_45_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_45_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_45_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_45_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_45_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_45_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_45_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_45_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_46_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_46_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_46_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_46_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_46_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_46_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_46_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_46_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_46_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_46_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_46_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_46_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_46_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_46_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_46_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_46_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_46_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_46_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_47_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_47_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_47_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_47_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_47_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_47_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_47_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_47_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_47_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_47_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_47_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_47_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_47_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_47_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_47_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_47_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_47_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_47_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_48_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_48_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_48_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_48_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_48_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_48_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_48_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_48_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_48_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_48_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_48_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_48_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_48_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_48_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_48_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_48_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_48_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_48_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_49_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_49_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_49_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_49_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_49_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_49_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_49_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_49_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_49_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_49_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_49_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_49_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_49_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_49_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_49_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_49_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_49_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_49_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_50_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_50_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_50_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_50_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_50_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_50_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_50_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_50_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_50_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_50_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_50_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_50_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_50_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_50_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_50_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_50_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_50_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_50_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_51_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_51_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_51_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_51_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_51_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_51_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_51_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_51_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_51_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_51_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_51_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_51_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_51_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_51_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_51_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_51_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_51_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_51_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_52_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_52_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_52_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_52_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_52_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_52_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_52_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_52_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_52_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_52_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_52_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_52_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_52_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_52_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_52_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_52_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_52_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_52_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_53_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_53_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_53_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_53_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_53_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_53_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_53_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_53_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_53_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_53_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_53_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_53_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_53_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_53_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_53_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_53_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_53_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_53_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_54_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_54_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_54_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_54_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_54_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_54_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_54_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_54_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_54_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_54_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_54_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_54_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_54_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_54_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_54_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_54_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_54_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_54_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_55_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_55_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_55_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_55_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_55_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_55_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_55_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_55_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_55_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_55_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_55_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_55_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_55_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_55_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_55_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_55_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_55_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_55_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_56_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_56_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_56_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_56_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_56_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_56_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_56_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_56_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_56_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_56_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_56_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_56_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_56_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_56_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_56_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_56_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_56_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_56_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_57_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_57_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_57_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_57_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_57_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_57_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_57_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_57_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_57_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_57_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_57_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_57_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_57_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_57_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_57_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_57_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_57_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_57_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_58_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_58_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_58_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_58_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_58_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_58_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_58_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_58_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_58_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_58_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_58_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_58_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_58_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_58_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_58_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_58_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_58_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_58_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_59_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_59_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_59_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_59_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_59_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_59_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_59_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_59_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_59_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_59_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_59_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_59_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_59_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_59_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_59_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_59_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_59_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_59_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_60_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_60_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_60_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_60_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_60_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_60_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_60_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_60_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_60_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_60_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_60_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_60_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_60_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_60_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_60_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_60_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_60_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_60_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_61_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_61_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_61_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_61_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_61_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_61_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_61_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_61_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_61_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_61_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_61_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_61_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_61_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_61_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_61_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_61_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_61_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_61_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_62_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_62_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_62_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_62_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_62_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_62_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_62_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_62_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_62_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_62_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_62_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_62_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_62_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_62_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_62_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_62_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_62_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_62_data_MPORT_3_addr_pipe_0;
  reg  inputDataBuffer_63_validBit [0:255]; // @[BP.scala 42:36]
  wire  inputDataBuffer_63_validBit_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_63_validBit_MPORT_3_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_63_validBit_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_63_validBit_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_63_validBit_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_63_validBit_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_63_validBit_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_63_validBit_MPORT_3_addr_pipe_0;
  reg [3:0] inputDataBuffer_63_data [0:255]; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_63_data_MPORT_3_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_63_data_MPORT_3_addr; // @[BP.scala 42:36]
  wire [3:0] inputDataBuffer_63_data_MPORT_data; // @[BP.scala 42:36]
  wire [7:0] inputDataBuffer_63_data_MPORT_addr; // @[BP.scala 42:36]
  wire  inputDataBuffer_63_data_MPORT_mask; // @[BP.scala 42:36]
  wire  inputDataBuffer_63_data_MPORT_en; // @[BP.scala 42:36]
  reg  inputDataBuffer_63_data_MPORT_3_en_pipe_0;
  reg [7:0] inputDataBuffer_63_data_MPORT_3_addr_pipe_0;
  wire  array_0_clock; // @[BP.scala 45:51]
  wire  array_0_reset; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_0_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_0_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_0_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_0_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_0_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_0_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_0_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_0_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_0_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_0_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_0_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_0_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_0_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_0_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_0_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_0_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_0_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_0_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_0_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_0_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_0_io_Addr_out; // @[BP.scala 45:51]
  wire  array_1_clock; // @[BP.scala 45:51]
  wire  array_1_reset; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_1_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_1_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_1_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_1_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_1_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_1_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_1_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_1_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_1_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_1_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_1_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_1_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_1_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_1_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_1_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_1_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_1_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_1_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_1_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_1_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_1_io_Addr_out; // @[BP.scala 45:51]
  wire  array_2_clock; // @[BP.scala 45:51]
  wire  array_2_reset; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_2_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_2_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_2_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_2_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_2_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_2_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_2_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_2_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_2_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_2_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_2_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_2_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_2_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_2_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_2_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_2_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_2_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_2_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_2_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_2_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_2_io_Addr_out; // @[BP.scala 45:51]
  wire  array_3_clock; // @[BP.scala 45:51]
  wire  array_3_reset; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_3_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_3_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_3_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_3_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_3_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_3_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_3_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_3_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_3_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_3_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_3_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_3_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_3_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_3_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_3_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_3_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_3_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_3_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_3_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_3_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_3_io_Addr_out; // @[BP.scala 45:51]
  wire  array_4_clock; // @[BP.scala 45:51]
  wire  array_4_reset; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_4_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_4_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_4_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_4_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_4_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_4_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_4_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_4_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_4_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_4_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_4_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_4_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_4_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_4_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_4_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_4_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_4_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_4_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_4_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_4_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_4_io_Addr_out; // @[BP.scala 45:51]
  wire  array_5_clock; // @[BP.scala 45:51]
  wire  array_5_reset; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_5_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_5_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_5_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_5_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_5_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_5_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_5_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_5_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_5_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_5_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_5_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_5_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_5_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_5_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_5_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_5_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_5_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_5_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_5_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_5_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_5_io_Addr_out; // @[BP.scala 45:51]
  wire  array_6_clock; // @[BP.scala 45:51]
  wire  array_6_reset; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_6_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_6_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_6_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_6_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_6_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_6_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_6_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_6_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_6_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_6_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_6_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_6_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_6_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_6_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_6_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_6_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_6_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_6_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_6_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_6_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_6_io_Addr_out; // @[BP.scala 45:51]
  wire  array_7_clock; // @[BP.scala 45:51]
  wire  array_7_reset; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_7_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_7_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_7_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_7_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_7_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_7_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_7_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_7_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_7_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_7_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_7_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_7_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_7_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_7_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_7_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_7_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_7_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_7_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_7_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_7_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_7_io_Addr_out; // @[BP.scala 45:51]
  wire  array_8_clock; // @[BP.scala 45:51]
  wire  array_8_reset; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_8_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_8_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_8_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_8_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_8_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_8_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_8_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_8_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_8_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_8_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_8_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_8_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_8_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_8_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_8_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_8_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_8_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_8_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_8_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_8_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_8_io_Addr_out; // @[BP.scala 45:51]
  wire  array_9_clock; // @[BP.scala 45:51]
  wire  array_9_reset; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_9_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_9_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_9_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_9_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_9_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_9_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_9_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_9_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_9_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_9_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_9_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_9_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_9_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_9_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_9_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_9_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_9_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_9_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_9_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_9_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_9_io_Addr_out; // @[BP.scala 45:51]
  wire  array_10_clock; // @[BP.scala 45:51]
  wire  array_10_reset; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_10_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_10_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_10_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_10_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_10_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_10_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_10_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_10_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_10_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_10_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_10_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_10_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_10_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_10_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_10_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_10_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_10_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_10_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_10_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_10_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_10_io_Addr_out; // @[BP.scala 45:51]
  wire  array_11_clock; // @[BP.scala 45:51]
  wire  array_11_reset; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_11_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_11_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_11_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_11_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_11_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_11_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_11_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_11_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_11_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_11_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_11_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_11_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_11_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_11_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_11_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_11_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_11_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_11_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_11_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_11_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_11_io_Addr_out; // @[BP.scala 45:51]
  wire  array_12_clock; // @[BP.scala 45:51]
  wire  array_12_reset; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_12_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_12_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_12_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_12_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_12_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_12_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_12_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_12_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_12_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_12_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_12_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_12_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_12_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_12_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_12_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_12_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_12_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_12_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_12_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_12_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_12_io_Addr_out; // @[BP.scala 45:51]
  wire  array_13_clock; // @[BP.scala 45:51]
  wire  array_13_reset; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_13_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_13_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_13_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_13_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_13_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_13_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_13_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_13_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_13_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_13_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_13_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_13_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_13_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_13_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_13_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_13_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_13_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_13_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_13_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_13_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_13_io_Addr_out; // @[BP.scala 45:51]
  wire  array_14_clock; // @[BP.scala 45:51]
  wire  array_14_reset; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_14_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_14_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_14_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_14_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_14_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_14_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_14_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_14_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_14_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_14_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_14_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_14_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_14_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_14_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_14_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_14_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_14_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_14_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_14_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_14_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_14_io_Addr_out; // @[BP.scala 45:51]
  wire  array_15_clock; // @[BP.scala 45:51]
  wire  array_15_reset; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_15_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_15_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_15_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_15_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_15_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_15_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_15_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_15_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_15_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_15_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_15_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_15_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_15_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_15_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_15_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_15_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_15_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_15_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_15_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_15_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_15_io_Addr_out; // @[BP.scala 45:51]
  wire  array_16_clock; // @[BP.scala 45:51]
  wire  array_16_reset; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_16_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_16_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_16_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_16_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_16_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_16_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_16_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_16_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_16_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_16_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_16_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_16_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_16_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_16_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_16_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_16_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_16_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_16_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_16_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_16_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_16_io_Addr_out; // @[BP.scala 45:51]
  wire  array_17_clock; // @[BP.scala 45:51]
  wire  array_17_reset; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_17_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_17_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_17_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_17_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_17_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_17_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_17_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_17_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_17_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_17_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_17_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_17_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_17_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_17_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_17_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_17_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_17_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_17_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_17_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_17_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_17_io_Addr_out; // @[BP.scala 45:51]
  wire  array_18_clock; // @[BP.scala 45:51]
  wire  array_18_reset; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_18_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_18_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_18_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_18_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_18_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_18_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_18_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_18_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_18_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_18_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_18_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_18_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_18_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_18_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_18_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_18_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_18_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_18_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_18_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_18_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_18_io_Addr_out; // @[BP.scala 45:51]
  wire  array_19_clock; // @[BP.scala 45:51]
  wire  array_19_reset; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_19_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_19_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_19_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_19_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_19_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_19_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_19_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_19_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_19_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_19_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_19_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_19_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_19_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_19_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_19_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_19_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_19_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_19_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_19_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_19_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_19_io_Addr_out; // @[BP.scala 45:51]
  wire  array_20_clock; // @[BP.scala 45:51]
  wire  array_20_reset; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_0_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_0_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_1_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_1_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_2_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_2_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_3_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_3_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_4_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_4_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_5_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_5_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_6_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_6_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_7_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_7_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_8_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_8_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_9_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_9_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_10_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_10_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_11_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_11_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_12_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_12_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_13_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_13_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_14_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_14_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_15_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_15_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_16_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_16_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_17_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_17_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_18_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_18_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_19_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_19_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_20_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_20_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_21_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_21_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_22_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_22_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_23_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_23_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_24_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_24_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_25_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_25_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_26_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_26_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_27_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_27_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_28_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_28_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_29_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_29_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_30_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_30_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_31_a; // @[BP.scala 45:51]
  wire  array_20_io_d_in_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_in_31_b; // @[BP.scala 45:51]
  wire  array_20_io_d_in_31_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_0_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_0_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_0_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_0_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_1_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_1_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_1_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_1_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_2_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_2_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_2_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_2_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_3_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_3_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_3_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_3_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_4_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_4_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_4_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_4_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_5_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_5_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_5_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_5_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_6_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_6_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_6_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_6_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_7_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_7_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_7_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_7_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_8_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_8_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_8_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_8_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_9_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_9_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_9_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_9_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_10_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_10_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_10_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_10_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_11_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_11_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_11_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_11_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_12_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_12_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_12_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_12_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_13_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_13_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_13_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_13_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_14_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_14_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_14_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_14_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_15_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_15_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_15_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_15_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_16_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_16_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_16_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_16_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_17_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_17_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_17_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_17_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_18_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_18_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_18_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_18_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_19_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_19_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_19_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_19_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_20_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_20_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_20_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_20_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_21_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_21_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_21_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_21_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_22_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_22_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_22_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_22_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_23_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_23_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_23_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_23_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_24_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_24_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_24_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_24_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_25_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_25_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_25_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_25_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_26_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_26_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_26_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_26_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_27_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_27_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_27_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_27_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_28_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_28_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_28_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_28_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_29_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_29_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_29_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_29_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_30_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_30_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_30_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_30_valid_b; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_31_a; // @[BP.scala 45:51]
  wire  array_20_io_d_out_31_valid_a; // @[BP.scala 45:51]
  wire [3:0] array_20_io_d_out_31_b; // @[BP.scala 45:51]
  wire  array_20_io_d_out_31_valid_b; // @[BP.scala 45:51]
  wire  array_20_io_wr_en_mem1; // @[BP.scala 45:51]
  wire  array_20_io_wr_en_mem2; // @[BP.scala 45:51]
  wire  array_20_io_wr_en_mem3; // @[BP.scala 45:51]
  wire  array_20_io_wr_en_mem4; // @[BP.scala 45:51]
  wire  array_20_io_wr_en_mem5; // @[BP.scala 45:51]
  wire  array_20_io_wr_en_mem6; // @[BP.scala 45:51]
  wire [287:0] array_20_io_wr_instr_mem1; // @[BP.scala 45:51]
  wire [127:0] array_20_io_wr_instr_mem2; // @[BP.scala 45:51]
  wire [127:0] array_20_io_wr_instr_mem3; // @[BP.scala 45:51]
  wire [127:0] array_20_io_wr_instr_mem4; // @[BP.scala 45:51]
  wire [127:0] array_20_io_wr_instr_mem5; // @[BP.scala 45:51]
  wire [127:0] array_20_io_wr_instr_mem6; // @[BP.scala 45:51]
  wire [7:0] array_20_io_PC1_in; // @[BP.scala 45:51]
  wire [7:0] array_20_io_PC6_out; // @[BP.scala 45:51]
  wire [7:0] array_20_io_Addr_in; // @[BP.scala 45:51]
  wire [7:0] array_20_io_Addr_out; // @[BP.scala 45:51]
  reg  outputDataBuffer_0_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_0_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_0_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_0_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_0_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_0_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_0_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_0_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_0_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_0_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_0_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_0_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_0_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_0_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_0_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_0_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_1_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_1_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_1_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_1_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_1_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_1_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_1_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_1_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_1_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_1_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_1_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_1_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_1_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_1_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_1_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_1_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_2_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_2_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_2_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_2_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_2_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_2_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_2_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_2_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_2_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_2_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_2_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_2_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_2_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_2_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_2_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_2_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_3_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_3_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_3_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_3_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_3_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_3_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_3_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_3_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_3_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_3_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_3_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_3_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_3_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_3_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_3_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_3_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_4_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_4_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_4_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_4_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_4_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_4_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_4_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_4_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_4_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_4_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_4_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_4_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_4_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_4_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_4_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_4_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_5_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_5_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_5_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_5_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_5_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_5_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_5_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_5_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_5_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_5_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_5_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_5_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_5_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_5_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_5_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_5_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_6_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_6_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_6_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_6_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_6_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_6_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_6_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_6_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_6_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_6_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_6_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_6_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_6_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_6_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_6_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_6_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_7_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_7_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_7_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_7_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_7_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_7_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_7_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_7_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_7_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_7_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_7_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_7_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_7_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_7_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_7_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_7_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_8_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_8_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_8_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_8_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_8_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_8_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_8_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_8_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_8_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_8_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_8_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_8_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_8_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_8_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_8_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_8_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_9_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_9_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_9_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_9_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_9_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_9_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_9_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_9_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_9_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_9_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_9_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_9_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_9_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_9_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_9_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_9_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_10_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_10_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_10_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_10_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_10_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_10_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_10_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_10_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_10_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_10_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_10_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_10_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_10_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_10_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_10_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_10_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_11_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_11_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_11_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_11_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_11_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_11_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_11_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_11_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_11_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_11_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_11_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_11_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_11_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_11_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_11_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_11_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_12_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_12_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_12_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_12_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_12_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_12_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_12_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_12_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_12_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_12_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_12_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_12_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_12_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_12_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_12_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_12_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_13_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_13_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_13_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_13_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_13_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_13_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_13_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_13_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_13_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_13_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_13_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_13_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_13_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_13_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_13_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_13_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_14_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_14_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_14_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_14_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_14_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_14_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_14_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_14_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_14_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_14_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_14_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_14_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_14_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_14_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_14_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_14_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_15_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_15_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_15_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_15_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_15_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_15_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_15_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_15_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_15_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_15_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_15_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_15_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_15_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_15_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_15_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_15_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_16_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_16_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_16_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_16_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_16_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_16_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_16_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_16_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_16_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_16_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_16_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_16_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_16_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_16_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_16_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_16_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_17_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_17_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_17_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_17_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_17_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_17_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_17_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_17_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_17_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_17_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_17_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_17_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_17_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_17_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_17_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_17_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_18_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_18_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_18_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_18_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_18_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_18_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_18_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_18_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_18_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_18_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_18_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_18_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_18_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_18_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_18_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_18_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_19_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_19_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_19_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_19_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_19_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_19_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_19_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_19_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_19_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_19_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_19_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_19_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_19_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_19_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_19_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_19_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_20_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_20_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_20_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_20_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_20_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_20_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_20_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_20_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_20_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_20_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_20_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_20_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_20_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_20_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_20_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_20_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_21_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_21_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_21_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_21_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_21_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_21_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_21_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_21_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_21_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_21_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_21_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_21_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_21_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_21_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_21_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_21_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_22_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_22_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_22_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_22_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_22_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_22_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_22_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_22_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_22_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_22_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_22_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_22_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_22_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_22_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_22_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_22_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_23_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_23_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_23_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_23_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_23_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_23_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_23_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_23_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_23_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_23_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_23_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_23_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_23_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_23_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_23_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_23_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_24_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_24_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_24_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_24_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_24_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_24_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_24_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_24_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_24_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_24_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_24_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_24_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_24_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_24_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_24_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_24_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_25_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_25_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_25_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_25_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_25_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_25_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_25_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_25_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_25_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_25_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_25_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_25_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_25_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_25_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_25_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_25_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_26_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_26_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_26_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_26_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_26_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_26_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_26_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_26_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_26_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_26_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_26_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_26_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_26_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_26_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_26_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_26_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_27_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_27_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_27_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_27_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_27_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_27_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_27_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_27_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_27_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_27_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_27_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_27_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_27_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_27_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_27_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_27_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_28_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_28_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_28_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_28_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_28_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_28_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_28_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_28_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_28_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_28_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_28_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_28_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_28_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_28_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_28_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_28_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_29_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_29_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_29_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_29_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_29_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_29_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_29_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_29_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_29_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_29_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_29_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_29_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_29_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_29_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_29_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_29_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_30_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_30_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_30_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_30_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_30_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_30_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_30_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_30_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_30_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_30_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_30_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_30_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_30_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_30_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_30_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_30_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_31_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_31_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_31_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_31_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_31_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_31_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_31_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_31_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_31_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_31_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_31_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_31_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_31_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_31_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_31_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_31_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_32_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_32_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_32_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_32_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_32_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_32_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_32_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_32_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_32_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_32_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_32_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_32_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_32_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_32_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_32_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_32_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_33_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_33_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_33_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_33_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_33_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_33_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_33_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_33_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_33_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_33_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_33_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_33_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_33_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_33_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_33_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_33_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_34_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_34_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_34_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_34_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_34_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_34_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_34_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_34_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_34_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_34_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_34_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_34_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_34_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_34_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_34_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_34_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_35_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_35_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_35_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_35_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_35_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_35_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_35_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_35_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_35_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_35_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_35_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_35_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_35_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_35_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_35_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_35_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_36_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_36_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_36_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_36_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_36_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_36_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_36_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_36_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_36_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_36_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_36_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_36_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_36_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_36_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_36_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_36_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_37_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_37_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_37_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_37_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_37_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_37_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_37_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_37_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_37_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_37_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_37_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_37_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_37_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_37_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_37_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_37_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_38_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_38_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_38_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_38_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_38_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_38_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_38_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_38_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_38_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_38_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_38_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_38_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_38_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_38_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_38_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_38_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_39_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_39_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_39_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_39_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_39_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_39_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_39_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_39_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_39_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_39_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_39_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_39_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_39_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_39_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_39_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_39_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_40_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_40_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_40_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_40_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_40_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_40_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_40_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_40_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_40_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_40_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_40_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_40_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_40_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_40_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_40_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_40_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_41_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_41_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_41_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_41_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_41_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_41_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_41_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_41_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_41_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_41_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_41_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_41_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_41_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_41_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_41_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_41_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_42_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_42_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_42_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_42_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_42_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_42_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_42_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_42_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_42_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_42_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_42_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_42_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_42_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_42_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_42_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_42_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_43_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_43_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_43_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_43_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_43_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_43_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_43_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_43_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_43_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_43_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_43_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_43_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_43_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_43_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_43_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_43_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_44_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_44_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_44_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_44_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_44_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_44_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_44_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_44_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_44_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_44_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_44_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_44_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_44_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_44_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_44_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_44_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_45_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_45_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_45_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_45_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_45_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_45_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_45_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_45_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_45_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_45_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_45_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_45_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_45_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_45_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_45_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_45_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_46_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_46_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_46_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_46_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_46_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_46_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_46_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_46_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_46_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_46_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_46_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_46_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_46_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_46_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_46_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_46_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_47_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_47_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_47_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_47_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_47_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_47_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_47_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_47_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_47_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_47_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_47_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_47_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_47_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_47_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_47_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_47_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_48_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_48_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_48_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_48_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_48_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_48_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_48_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_48_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_48_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_48_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_48_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_48_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_48_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_48_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_48_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_48_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_49_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_49_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_49_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_49_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_49_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_49_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_49_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_49_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_49_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_49_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_49_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_49_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_49_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_49_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_49_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_49_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_50_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_50_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_50_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_50_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_50_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_50_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_50_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_50_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_50_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_50_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_50_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_50_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_50_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_50_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_50_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_50_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_51_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_51_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_51_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_51_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_51_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_51_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_51_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_51_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_51_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_51_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_51_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_51_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_51_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_51_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_51_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_51_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_52_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_52_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_52_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_52_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_52_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_52_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_52_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_52_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_52_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_52_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_52_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_52_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_52_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_52_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_52_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_52_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_53_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_53_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_53_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_53_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_53_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_53_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_53_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_53_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_53_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_53_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_53_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_53_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_53_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_53_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_53_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_53_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_54_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_54_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_54_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_54_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_54_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_54_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_54_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_54_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_54_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_54_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_54_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_54_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_54_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_54_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_54_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_54_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_55_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_55_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_55_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_55_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_55_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_55_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_55_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_55_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_55_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_55_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_55_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_55_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_55_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_55_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_55_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_55_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_56_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_56_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_56_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_56_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_56_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_56_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_56_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_56_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_56_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_56_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_56_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_56_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_56_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_56_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_56_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_56_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_57_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_57_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_57_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_57_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_57_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_57_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_57_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_57_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_57_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_57_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_57_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_57_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_57_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_57_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_57_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_57_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_58_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_58_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_58_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_58_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_58_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_58_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_58_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_58_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_58_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_58_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_58_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_58_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_58_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_58_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_58_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_58_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_59_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_59_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_59_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_59_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_59_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_59_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_59_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_59_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_59_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_59_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_59_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_59_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_59_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_59_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_59_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_59_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_60_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_60_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_60_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_60_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_60_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_60_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_60_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_60_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_60_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_60_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_60_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_60_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_60_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_60_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_60_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_60_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_61_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_61_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_61_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_61_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_61_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_61_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_61_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_61_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_61_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_61_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_61_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_61_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_61_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_61_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_61_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_61_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_62_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_62_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_62_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_62_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_62_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_62_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_62_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_62_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_62_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_62_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_62_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_62_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_62_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_62_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_62_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_62_data_MPORT_2_addr_pipe_0;
  reg  outputDataBuffer_63_validBit [0:255]; // @[BP.scala 47:37]
  wire  outputDataBuffer_63_validBit_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_63_validBit_MPORT_2_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_63_validBit_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_63_validBit_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_63_validBit_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_63_validBit_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_63_validBit_MPORT_2_addr_pipe_0;
  reg [3:0] outputDataBuffer_63_data [0:255]; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_63_data_MPORT_2_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_63_data_MPORT_2_addr; // @[BP.scala 47:37]
  wire [3:0] outputDataBuffer_63_data_MPORT_4_data; // @[BP.scala 47:37]
  wire [7:0] outputDataBuffer_63_data_MPORT_4_addr; // @[BP.scala 47:37]
  wire  outputDataBuffer_63_data_MPORT_4_mask; // @[BP.scala 47:37]
  wire  outputDataBuffer_63_data_MPORT_4_en; // @[BP.scala 47:37]
  reg [7:0] outputDataBuffer_63_data_MPORT_2_addr_pipe_0;
  reg [7:0] wr_Addr_inBuf; // @[BP.scala 50:30]
  wire [7:0] _wr_Addr_inBuf_T_1 = wr_Addr_inBuf + 8'h1; // @[BP.scala 61:36]
  reg [7:0] rd_Addr_inBuf; // @[BP.scala 91:30]
  reg  rd_D_inBuf_0_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_0_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_1_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_1_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_2_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_2_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_3_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_3_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_4_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_4_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_5_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_5_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_6_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_6_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_7_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_7_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_8_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_8_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_9_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_9_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_10_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_10_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_11_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_11_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_12_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_12_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_13_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_13_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_14_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_14_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_15_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_15_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_16_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_16_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_17_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_17_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_18_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_18_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_19_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_19_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_20_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_20_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_21_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_21_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_22_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_22_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_23_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_23_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_24_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_24_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_25_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_25_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_26_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_26_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_27_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_27_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_28_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_28_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_29_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_29_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_30_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_30_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_31_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_31_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_32_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_32_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_33_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_33_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_34_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_34_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_35_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_35_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_36_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_36_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_37_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_37_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_38_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_38_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_39_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_39_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_40_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_40_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_41_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_41_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_42_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_42_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_43_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_43_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_44_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_44_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_45_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_45_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_46_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_46_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_47_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_47_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_48_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_48_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_49_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_49_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_50_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_50_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_51_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_51_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_52_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_52_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_53_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_53_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_54_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_54_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_55_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_55_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_56_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_56_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_57_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_57_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_58_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_58_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_59_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_59_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_60_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_60_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_61_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_61_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_62_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_62_data; // @[BP.scala 93:23]
  reg  rd_D_inBuf_63_validBit; // @[BP.scala 93:23]
  reg [3:0] rd_D_inBuf_63_data; // @[BP.scala 93:23]
  wire [7:0] _rd_Addr_inBuf_T_1 = rd_Addr_inBuf + 8'h1; // @[BP.scala 101:36]
  reg [7:0] wr_Addr_outBuf; // @[BP.scala 114:31]
  reg  wr_D_outBuf_0_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_0_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_1_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_1_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_2_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_2_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_3_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_3_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_4_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_4_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_5_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_5_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_6_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_6_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_7_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_7_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_8_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_8_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_9_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_9_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_10_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_10_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_11_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_11_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_12_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_12_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_13_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_13_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_14_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_14_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_15_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_15_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_16_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_16_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_17_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_17_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_18_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_18_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_19_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_19_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_20_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_20_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_21_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_21_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_22_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_22_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_23_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_23_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_24_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_24_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_25_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_25_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_26_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_26_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_27_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_27_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_28_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_28_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_29_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_29_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_30_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_30_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_31_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_31_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_32_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_32_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_33_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_33_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_34_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_34_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_35_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_35_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_36_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_36_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_37_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_37_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_38_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_38_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_39_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_39_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_40_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_40_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_41_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_41_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_42_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_42_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_43_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_43_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_44_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_44_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_45_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_45_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_46_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_46_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_47_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_47_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_48_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_48_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_49_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_49_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_50_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_50_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_51_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_51_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_52_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_52_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_53_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_53_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_54_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_54_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_55_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_55_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_56_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_56_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_57_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_57_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_58_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_58_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_59_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_59_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_60_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_60_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_61_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_61_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_62_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_62_data; // @[BP.scala 117:24]
  reg  wr_D_outBuf_63_validBit; // @[BP.scala 117:24]
  reg [3:0] wr_D_outBuf_63_data; // @[BP.scala 117:24]
  reg [7:0] PCBegin; // @[BP.scala 287:24]
  reg [7:0] AddrBegin; // @[BP.scala 288:26]
  wire [7:0] _PCBegin_T_1 = PCBegin + 8'h1; // @[BP.scala 295:24]
  wire [7:0] _AddrBegin_T_1 = AddrBegin + 8'h1; // @[BP.scala 299:28]
  wire [7:0] Addr_out = array_20_io_Addr_out; // @[BP.scala 120:22 BP.scala 344:12]
  BuildingBlockNew array_0 ( // @[BP.scala 45:51]
    .clock(array_0_clock),
    .reset(array_0_reset),
    .io_d_in_0_a(array_0_io_d_in_0_a),
    .io_d_in_0_valid_a(array_0_io_d_in_0_valid_a),
    .io_d_in_0_b(array_0_io_d_in_0_b),
    .io_d_in_0_valid_b(array_0_io_d_in_0_valid_b),
    .io_d_in_1_a(array_0_io_d_in_1_a),
    .io_d_in_1_valid_a(array_0_io_d_in_1_valid_a),
    .io_d_in_1_b(array_0_io_d_in_1_b),
    .io_d_in_1_valid_b(array_0_io_d_in_1_valid_b),
    .io_d_in_2_a(array_0_io_d_in_2_a),
    .io_d_in_2_valid_a(array_0_io_d_in_2_valid_a),
    .io_d_in_2_b(array_0_io_d_in_2_b),
    .io_d_in_2_valid_b(array_0_io_d_in_2_valid_b),
    .io_d_in_3_a(array_0_io_d_in_3_a),
    .io_d_in_3_valid_a(array_0_io_d_in_3_valid_a),
    .io_d_in_3_b(array_0_io_d_in_3_b),
    .io_d_in_3_valid_b(array_0_io_d_in_3_valid_b),
    .io_d_in_4_a(array_0_io_d_in_4_a),
    .io_d_in_4_valid_a(array_0_io_d_in_4_valid_a),
    .io_d_in_4_b(array_0_io_d_in_4_b),
    .io_d_in_4_valid_b(array_0_io_d_in_4_valid_b),
    .io_d_in_5_a(array_0_io_d_in_5_a),
    .io_d_in_5_valid_a(array_0_io_d_in_5_valid_a),
    .io_d_in_5_b(array_0_io_d_in_5_b),
    .io_d_in_5_valid_b(array_0_io_d_in_5_valid_b),
    .io_d_in_6_a(array_0_io_d_in_6_a),
    .io_d_in_6_valid_a(array_0_io_d_in_6_valid_a),
    .io_d_in_6_b(array_0_io_d_in_6_b),
    .io_d_in_6_valid_b(array_0_io_d_in_6_valid_b),
    .io_d_in_7_a(array_0_io_d_in_7_a),
    .io_d_in_7_valid_a(array_0_io_d_in_7_valid_a),
    .io_d_in_7_b(array_0_io_d_in_7_b),
    .io_d_in_7_valid_b(array_0_io_d_in_7_valid_b),
    .io_d_in_8_a(array_0_io_d_in_8_a),
    .io_d_in_8_valid_a(array_0_io_d_in_8_valid_a),
    .io_d_in_8_b(array_0_io_d_in_8_b),
    .io_d_in_8_valid_b(array_0_io_d_in_8_valid_b),
    .io_d_in_9_a(array_0_io_d_in_9_a),
    .io_d_in_9_valid_a(array_0_io_d_in_9_valid_a),
    .io_d_in_9_b(array_0_io_d_in_9_b),
    .io_d_in_9_valid_b(array_0_io_d_in_9_valid_b),
    .io_d_in_10_a(array_0_io_d_in_10_a),
    .io_d_in_10_valid_a(array_0_io_d_in_10_valid_a),
    .io_d_in_10_b(array_0_io_d_in_10_b),
    .io_d_in_10_valid_b(array_0_io_d_in_10_valid_b),
    .io_d_in_11_a(array_0_io_d_in_11_a),
    .io_d_in_11_valid_a(array_0_io_d_in_11_valid_a),
    .io_d_in_11_b(array_0_io_d_in_11_b),
    .io_d_in_11_valid_b(array_0_io_d_in_11_valid_b),
    .io_d_in_12_a(array_0_io_d_in_12_a),
    .io_d_in_12_valid_a(array_0_io_d_in_12_valid_a),
    .io_d_in_12_b(array_0_io_d_in_12_b),
    .io_d_in_12_valid_b(array_0_io_d_in_12_valid_b),
    .io_d_in_13_a(array_0_io_d_in_13_a),
    .io_d_in_13_valid_a(array_0_io_d_in_13_valid_a),
    .io_d_in_13_b(array_0_io_d_in_13_b),
    .io_d_in_13_valid_b(array_0_io_d_in_13_valid_b),
    .io_d_in_14_a(array_0_io_d_in_14_a),
    .io_d_in_14_valid_a(array_0_io_d_in_14_valid_a),
    .io_d_in_14_b(array_0_io_d_in_14_b),
    .io_d_in_14_valid_b(array_0_io_d_in_14_valid_b),
    .io_d_in_15_a(array_0_io_d_in_15_a),
    .io_d_in_15_valid_a(array_0_io_d_in_15_valid_a),
    .io_d_in_15_b(array_0_io_d_in_15_b),
    .io_d_in_15_valid_b(array_0_io_d_in_15_valid_b),
    .io_d_in_16_a(array_0_io_d_in_16_a),
    .io_d_in_16_valid_a(array_0_io_d_in_16_valid_a),
    .io_d_in_16_b(array_0_io_d_in_16_b),
    .io_d_in_16_valid_b(array_0_io_d_in_16_valid_b),
    .io_d_in_17_a(array_0_io_d_in_17_a),
    .io_d_in_17_valid_a(array_0_io_d_in_17_valid_a),
    .io_d_in_17_b(array_0_io_d_in_17_b),
    .io_d_in_17_valid_b(array_0_io_d_in_17_valid_b),
    .io_d_in_18_a(array_0_io_d_in_18_a),
    .io_d_in_18_valid_a(array_0_io_d_in_18_valid_a),
    .io_d_in_18_b(array_0_io_d_in_18_b),
    .io_d_in_18_valid_b(array_0_io_d_in_18_valid_b),
    .io_d_in_19_a(array_0_io_d_in_19_a),
    .io_d_in_19_valid_a(array_0_io_d_in_19_valid_a),
    .io_d_in_19_b(array_0_io_d_in_19_b),
    .io_d_in_19_valid_b(array_0_io_d_in_19_valid_b),
    .io_d_in_20_a(array_0_io_d_in_20_a),
    .io_d_in_20_valid_a(array_0_io_d_in_20_valid_a),
    .io_d_in_20_b(array_0_io_d_in_20_b),
    .io_d_in_20_valid_b(array_0_io_d_in_20_valid_b),
    .io_d_in_21_a(array_0_io_d_in_21_a),
    .io_d_in_21_valid_a(array_0_io_d_in_21_valid_a),
    .io_d_in_21_b(array_0_io_d_in_21_b),
    .io_d_in_21_valid_b(array_0_io_d_in_21_valid_b),
    .io_d_in_22_a(array_0_io_d_in_22_a),
    .io_d_in_22_valid_a(array_0_io_d_in_22_valid_a),
    .io_d_in_22_b(array_0_io_d_in_22_b),
    .io_d_in_22_valid_b(array_0_io_d_in_22_valid_b),
    .io_d_in_23_a(array_0_io_d_in_23_a),
    .io_d_in_23_valid_a(array_0_io_d_in_23_valid_a),
    .io_d_in_23_b(array_0_io_d_in_23_b),
    .io_d_in_23_valid_b(array_0_io_d_in_23_valid_b),
    .io_d_in_24_a(array_0_io_d_in_24_a),
    .io_d_in_24_valid_a(array_0_io_d_in_24_valid_a),
    .io_d_in_24_b(array_0_io_d_in_24_b),
    .io_d_in_24_valid_b(array_0_io_d_in_24_valid_b),
    .io_d_in_25_a(array_0_io_d_in_25_a),
    .io_d_in_25_valid_a(array_0_io_d_in_25_valid_a),
    .io_d_in_25_b(array_0_io_d_in_25_b),
    .io_d_in_25_valid_b(array_0_io_d_in_25_valid_b),
    .io_d_in_26_a(array_0_io_d_in_26_a),
    .io_d_in_26_valid_a(array_0_io_d_in_26_valid_a),
    .io_d_in_26_b(array_0_io_d_in_26_b),
    .io_d_in_26_valid_b(array_0_io_d_in_26_valid_b),
    .io_d_in_27_a(array_0_io_d_in_27_a),
    .io_d_in_27_valid_a(array_0_io_d_in_27_valid_a),
    .io_d_in_27_b(array_0_io_d_in_27_b),
    .io_d_in_27_valid_b(array_0_io_d_in_27_valid_b),
    .io_d_in_28_a(array_0_io_d_in_28_a),
    .io_d_in_28_valid_a(array_0_io_d_in_28_valid_a),
    .io_d_in_28_b(array_0_io_d_in_28_b),
    .io_d_in_28_valid_b(array_0_io_d_in_28_valid_b),
    .io_d_in_29_a(array_0_io_d_in_29_a),
    .io_d_in_29_valid_a(array_0_io_d_in_29_valid_a),
    .io_d_in_29_b(array_0_io_d_in_29_b),
    .io_d_in_29_valid_b(array_0_io_d_in_29_valid_b),
    .io_d_in_30_a(array_0_io_d_in_30_a),
    .io_d_in_30_valid_a(array_0_io_d_in_30_valid_a),
    .io_d_in_30_b(array_0_io_d_in_30_b),
    .io_d_in_30_valid_b(array_0_io_d_in_30_valid_b),
    .io_d_in_31_a(array_0_io_d_in_31_a),
    .io_d_in_31_valid_a(array_0_io_d_in_31_valid_a),
    .io_d_in_31_b(array_0_io_d_in_31_b),
    .io_d_in_31_valid_b(array_0_io_d_in_31_valid_b),
    .io_d_out_0_a(array_0_io_d_out_0_a),
    .io_d_out_0_valid_a(array_0_io_d_out_0_valid_a),
    .io_d_out_0_b(array_0_io_d_out_0_b),
    .io_d_out_0_valid_b(array_0_io_d_out_0_valid_b),
    .io_d_out_1_a(array_0_io_d_out_1_a),
    .io_d_out_1_valid_a(array_0_io_d_out_1_valid_a),
    .io_d_out_1_b(array_0_io_d_out_1_b),
    .io_d_out_1_valid_b(array_0_io_d_out_1_valid_b),
    .io_d_out_2_a(array_0_io_d_out_2_a),
    .io_d_out_2_valid_a(array_0_io_d_out_2_valid_a),
    .io_d_out_2_b(array_0_io_d_out_2_b),
    .io_d_out_2_valid_b(array_0_io_d_out_2_valid_b),
    .io_d_out_3_a(array_0_io_d_out_3_a),
    .io_d_out_3_valid_a(array_0_io_d_out_3_valid_a),
    .io_d_out_3_b(array_0_io_d_out_3_b),
    .io_d_out_3_valid_b(array_0_io_d_out_3_valid_b),
    .io_d_out_4_a(array_0_io_d_out_4_a),
    .io_d_out_4_valid_a(array_0_io_d_out_4_valid_a),
    .io_d_out_4_b(array_0_io_d_out_4_b),
    .io_d_out_4_valid_b(array_0_io_d_out_4_valid_b),
    .io_d_out_5_a(array_0_io_d_out_5_a),
    .io_d_out_5_valid_a(array_0_io_d_out_5_valid_a),
    .io_d_out_5_b(array_0_io_d_out_5_b),
    .io_d_out_5_valid_b(array_0_io_d_out_5_valid_b),
    .io_d_out_6_a(array_0_io_d_out_6_a),
    .io_d_out_6_valid_a(array_0_io_d_out_6_valid_a),
    .io_d_out_6_b(array_0_io_d_out_6_b),
    .io_d_out_6_valid_b(array_0_io_d_out_6_valid_b),
    .io_d_out_7_a(array_0_io_d_out_7_a),
    .io_d_out_7_valid_a(array_0_io_d_out_7_valid_a),
    .io_d_out_7_b(array_0_io_d_out_7_b),
    .io_d_out_7_valid_b(array_0_io_d_out_7_valid_b),
    .io_d_out_8_a(array_0_io_d_out_8_a),
    .io_d_out_8_valid_a(array_0_io_d_out_8_valid_a),
    .io_d_out_8_b(array_0_io_d_out_8_b),
    .io_d_out_8_valid_b(array_0_io_d_out_8_valid_b),
    .io_d_out_9_a(array_0_io_d_out_9_a),
    .io_d_out_9_valid_a(array_0_io_d_out_9_valid_a),
    .io_d_out_9_b(array_0_io_d_out_9_b),
    .io_d_out_9_valid_b(array_0_io_d_out_9_valid_b),
    .io_d_out_10_a(array_0_io_d_out_10_a),
    .io_d_out_10_valid_a(array_0_io_d_out_10_valid_a),
    .io_d_out_10_b(array_0_io_d_out_10_b),
    .io_d_out_10_valid_b(array_0_io_d_out_10_valid_b),
    .io_d_out_11_a(array_0_io_d_out_11_a),
    .io_d_out_11_valid_a(array_0_io_d_out_11_valid_a),
    .io_d_out_11_b(array_0_io_d_out_11_b),
    .io_d_out_11_valid_b(array_0_io_d_out_11_valid_b),
    .io_d_out_12_a(array_0_io_d_out_12_a),
    .io_d_out_12_valid_a(array_0_io_d_out_12_valid_a),
    .io_d_out_12_b(array_0_io_d_out_12_b),
    .io_d_out_12_valid_b(array_0_io_d_out_12_valid_b),
    .io_d_out_13_a(array_0_io_d_out_13_a),
    .io_d_out_13_valid_a(array_0_io_d_out_13_valid_a),
    .io_d_out_13_b(array_0_io_d_out_13_b),
    .io_d_out_13_valid_b(array_0_io_d_out_13_valid_b),
    .io_d_out_14_a(array_0_io_d_out_14_a),
    .io_d_out_14_valid_a(array_0_io_d_out_14_valid_a),
    .io_d_out_14_b(array_0_io_d_out_14_b),
    .io_d_out_14_valid_b(array_0_io_d_out_14_valid_b),
    .io_d_out_15_a(array_0_io_d_out_15_a),
    .io_d_out_15_valid_a(array_0_io_d_out_15_valid_a),
    .io_d_out_15_b(array_0_io_d_out_15_b),
    .io_d_out_15_valid_b(array_0_io_d_out_15_valid_b),
    .io_d_out_16_a(array_0_io_d_out_16_a),
    .io_d_out_16_valid_a(array_0_io_d_out_16_valid_a),
    .io_d_out_16_b(array_0_io_d_out_16_b),
    .io_d_out_16_valid_b(array_0_io_d_out_16_valid_b),
    .io_d_out_17_a(array_0_io_d_out_17_a),
    .io_d_out_17_valid_a(array_0_io_d_out_17_valid_a),
    .io_d_out_17_b(array_0_io_d_out_17_b),
    .io_d_out_17_valid_b(array_0_io_d_out_17_valid_b),
    .io_d_out_18_a(array_0_io_d_out_18_a),
    .io_d_out_18_valid_a(array_0_io_d_out_18_valid_a),
    .io_d_out_18_b(array_0_io_d_out_18_b),
    .io_d_out_18_valid_b(array_0_io_d_out_18_valid_b),
    .io_d_out_19_a(array_0_io_d_out_19_a),
    .io_d_out_19_valid_a(array_0_io_d_out_19_valid_a),
    .io_d_out_19_b(array_0_io_d_out_19_b),
    .io_d_out_19_valid_b(array_0_io_d_out_19_valid_b),
    .io_d_out_20_a(array_0_io_d_out_20_a),
    .io_d_out_20_valid_a(array_0_io_d_out_20_valid_a),
    .io_d_out_20_b(array_0_io_d_out_20_b),
    .io_d_out_20_valid_b(array_0_io_d_out_20_valid_b),
    .io_d_out_21_a(array_0_io_d_out_21_a),
    .io_d_out_21_valid_a(array_0_io_d_out_21_valid_a),
    .io_d_out_21_b(array_0_io_d_out_21_b),
    .io_d_out_21_valid_b(array_0_io_d_out_21_valid_b),
    .io_d_out_22_a(array_0_io_d_out_22_a),
    .io_d_out_22_valid_a(array_0_io_d_out_22_valid_a),
    .io_d_out_22_b(array_0_io_d_out_22_b),
    .io_d_out_22_valid_b(array_0_io_d_out_22_valid_b),
    .io_d_out_23_a(array_0_io_d_out_23_a),
    .io_d_out_23_valid_a(array_0_io_d_out_23_valid_a),
    .io_d_out_23_b(array_0_io_d_out_23_b),
    .io_d_out_23_valid_b(array_0_io_d_out_23_valid_b),
    .io_d_out_24_a(array_0_io_d_out_24_a),
    .io_d_out_24_valid_a(array_0_io_d_out_24_valid_a),
    .io_d_out_24_b(array_0_io_d_out_24_b),
    .io_d_out_24_valid_b(array_0_io_d_out_24_valid_b),
    .io_d_out_25_a(array_0_io_d_out_25_a),
    .io_d_out_25_valid_a(array_0_io_d_out_25_valid_a),
    .io_d_out_25_b(array_0_io_d_out_25_b),
    .io_d_out_25_valid_b(array_0_io_d_out_25_valid_b),
    .io_d_out_26_a(array_0_io_d_out_26_a),
    .io_d_out_26_valid_a(array_0_io_d_out_26_valid_a),
    .io_d_out_26_b(array_0_io_d_out_26_b),
    .io_d_out_26_valid_b(array_0_io_d_out_26_valid_b),
    .io_d_out_27_a(array_0_io_d_out_27_a),
    .io_d_out_27_valid_a(array_0_io_d_out_27_valid_a),
    .io_d_out_27_b(array_0_io_d_out_27_b),
    .io_d_out_27_valid_b(array_0_io_d_out_27_valid_b),
    .io_d_out_28_a(array_0_io_d_out_28_a),
    .io_d_out_28_valid_a(array_0_io_d_out_28_valid_a),
    .io_d_out_28_b(array_0_io_d_out_28_b),
    .io_d_out_28_valid_b(array_0_io_d_out_28_valid_b),
    .io_d_out_29_a(array_0_io_d_out_29_a),
    .io_d_out_29_valid_a(array_0_io_d_out_29_valid_a),
    .io_d_out_29_b(array_0_io_d_out_29_b),
    .io_d_out_29_valid_b(array_0_io_d_out_29_valid_b),
    .io_d_out_30_a(array_0_io_d_out_30_a),
    .io_d_out_30_valid_a(array_0_io_d_out_30_valid_a),
    .io_d_out_30_b(array_0_io_d_out_30_b),
    .io_d_out_30_valid_b(array_0_io_d_out_30_valid_b),
    .io_d_out_31_a(array_0_io_d_out_31_a),
    .io_d_out_31_valid_a(array_0_io_d_out_31_valid_a),
    .io_d_out_31_b(array_0_io_d_out_31_b),
    .io_d_out_31_valid_b(array_0_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_0_io_wr_en_mem1),
    .io_wr_en_mem2(array_0_io_wr_en_mem2),
    .io_wr_en_mem3(array_0_io_wr_en_mem3),
    .io_wr_en_mem4(array_0_io_wr_en_mem4),
    .io_wr_en_mem5(array_0_io_wr_en_mem5),
    .io_wr_en_mem6(array_0_io_wr_en_mem6),
    .io_wr_instr_mem1(array_0_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_0_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_0_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_0_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_0_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_0_io_wr_instr_mem6),
    .io_PC1_in(array_0_io_PC1_in),
    .io_PC6_out(array_0_io_PC6_out),
    .io_Addr_in(array_0_io_Addr_in),
    .io_Addr_out(array_0_io_Addr_out)
  );
  BuildingBlockNew array_1 ( // @[BP.scala 45:51]
    .clock(array_1_clock),
    .reset(array_1_reset),
    .io_d_in_0_a(array_1_io_d_in_0_a),
    .io_d_in_0_valid_a(array_1_io_d_in_0_valid_a),
    .io_d_in_0_b(array_1_io_d_in_0_b),
    .io_d_in_0_valid_b(array_1_io_d_in_0_valid_b),
    .io_d_in_1_a(array_1_io_d_in_1_a),
    .io_d_in_1_valid_a(array_1_io_d_in_1_valid_a),
    .io_d_in_1_b(array_1_io_d_in_1_b),
    .io_d_in_1_valid_b(array_1_io_d_in_1_valid_b),
    .io_d_in_2_a(array_1_io_d_in_2_a),
    .io_d_in_2_valid_a(array_1_io_d_in_2_valid_a),
    .io_d_in_2_b(array_1_io_d_in_2_b),
    .io_d_in_2_valid_b(array_1_io_d_in_2_valid_b),
    .io_d_in_3_a(array_1_io_d_in_3_a),
    .io_d_in_3_valid_a(array_1_io_d_in_3_valid_a),
    .io_d_in_3_b(array_1_io_d_in_3_b),
    .io_d_in_3_valid_b(array_1_io_d_in_3_valid_b),
    .io_d_in_4_a(array_1_io_d_in_4_a),
    .io_d_in_4_valid_a(array_1_io_d_in_4_valid_a),
    .io_d_in_4_b(array_1_io_d_in_4_b),
    .io_d_in_4_valid_b(array_1_io_d_in_4_valid_b),
    .io_d_in_5_a(array_1_io_d_in_5_a),
    .io_d_in_5_valid_a(array_1_io_d_in_5_valid_a),
    .io_d_in_5_b(array_1_io_d_in_5_b),
    .io_d_in_5_valid_b(array_1_io_d_in_5_valid_b),
    .io_d_in_6_a(array_1_io_d_in_6_a),
    .io_d_in_6_valid_a(array_1_io_d_in_6_valid_a),
    .io_d_in_6_b(array_1_io_d_in_6_b),
    .io_d_in_6_valid_b(array_1_io_d_in_6_valid_b),
    .io_d_in_7_a(array_1_io_d_in_7_a),
    .io_d_in_7_valid_a(array_1_io_d_in_7_valid_a),
    .io_d_in_7_b(array_1_io_d_in_7_b),
    .io_d_in_7_valid_b(array_1_io_d_in_7_valid_b),
    .io_d_in_8_a(array_1_io_d_in_8_a),
    .io_d_in_8_valid_a(array_1_io_d_in_8_valid_a),
    .io_d_in_8_b(array_1_io_d_in_8_b),
    .io_d_in_8_valid_b(array_1_io_d_in_8_valid_b),
    .io_d_in_9_a(array_1_io_d_in_9_a),
    .io_d_in_9_valid_a(array_1_io_d_in_9_valid_a),
    .io_d_in_9_b(array_1_io_d_in_9_b),
    .io_d_in_9_valid_b(array_1_io_d_in_9_valid_b),
    .io_d_in_10_a(array_1_io_d_in_10_a),
    .io_d_in_10_valid_a(array_1_io_d_in_10_valid_a),
    .io_d_in_10_b(array_1_io_d_in_10_b),
    .io_d_in_10_valid_b(array_1_io_d_in_10_valid_b),
    .io_d_in_11_a(array_1_io_d_in_11_a),
    .io_d_in_11_valid_a(array_1_io_d_in_11_valid_a),
    .io_d_in_11_b(array_1_io_d_in_11_b),
    .io_d_in_11_valid_b(array_1_io_d_in_11_valid_b),
    .io_d_in_12_a(array_1_io_d_in_12_a),
    .io_d_in_12_valid_a(array_1_io_d_in_12_valid_a),
    .io_d_in_12_b(array_1_io_d_in_12_b),
    .io_d_in_12_valid_b(array_1_io_d_in_12_valid_b),
    .io_d_in_13_a(array_1_io_d_in_13_a),
    .io_d_in_13_valid_a(array_1_io_d_in_13_valid_a),
    .io_d_in_13_b(array_1_io_d_in_13_b),
    .io_d_in_13_valid_b(array_1_io_d_in_13_valid_b),
    .io_d_in_14_a(array_1_io_d_in_14_a),
    .io_d_in_14_valid_a(array_1_io_d_in_14_valid_a),
    .io_d_in_14_b(array_1_io_d_in_14_b),
    .io_d_in_14_valid_b(array_1_io_d_in_14_valid_b),
    .io_d_in_15_a(array_1_io_d_in_15_a),
    .io_d_in_15_valid_a(array_1_io_d_in_15_valid_a),
    .io_d_in_15_b(array_1_io_d_in_15_b),
    .io_d_in_15_valid_b(array_1_io_d_in_15_valid_b),
    .io_d_in_16_a(array_1_io_d_in_16_a),
    .io_d_in_16_valid_a(array_1_io_d_in_16_valid_a),
    .io_d_in_16_b(array_1_io_d_in_16_b),
    .io_d_in_16_valid_b(array_1_io_d_in_16_valid_b),
    .io_d_in_17_a(array_1_io_d_in_17_a),
    .io_d_in_17_valid_a(array_1_io_d_in_17_valid_a),
    .io_d_in_17_b(array_1_io_d_in_17_b),
    .io_d_in_17_valid_b(array_1_io_d_in_17_valid_b),
    .io_d_in_18_a(array_1_io_d_in_18_a),
    .io_d_in_18_valid_a(array_1_io_d_in_18_valid_a),
    .io_d_in_18_b(array_1_io_d_in_18_b),
    .io_d_in_18_valid_b(array_1_io_d_in_18_valid_b),
    .io_d_in_19_a(array_1_io_d_in_19_a),
    .io_d_in_19_valid_a(array_1_io_d_in_19_valid_a),
    .io_d_in_19_b(array_1_io_d_in_19_b),
    .io_d_in_19_valid_b(array_1_io_d_in_19_valid_b),
    .io_d_in_20_a(array_1_io_d_in_20_a),
    .io_d_in_20_valid_a(array_1_io_d_in_20_valid_a),
    .io_d_in_20_b(array_1_io_d_in_20_b),
    .io_d_in_20_valid_b(array_1_io_d_in_20_valid_b),
    .io_d_in_21_a(array_1_io_d_in_21_a),
    .io_d_in_21_valid_a(array_1_io_d_in_21_valid_a),
    .io_d_in_21_b(array_1_io_d_in_21_b),
    .io_d_in_21_valid_b(array_1_io_d_in_21_valid_b),
    .io_d_in_22_a(array_1_io_d_in_22_a),
    .io_d_in_22_valid_a(array_1_io_d_in_22_valid_a),
    .io_d_in_22_b(array_1_io_d_in_22_b),
    .io_d_in_22_valid_b(array_1_io_d_in_22_valid_b),
    .io_d_in_23_a(array_1_io_d_in_23_a),
    .io_d_in_23_valid_a(array_1_io_d_in_23_valid_a),
    .io_d_in_23_b(array_1_io_d_in_23_b),
    .io_d_in_23_valid_b(array_1_io_d_in_23_valid_b),
    .io_d_in_24_a(array_1_io_d_in_24_a),
    .io_d_in_24_valid_a(array_1_io_d_in_24_valid_a),
    .io_d_in_24_b(array_1_io_d_in_24_b),
    .io_d_in_24_valid_b(array_1_io_d_in_24_valid_b),
    .io_d_in_25_a(array_1_io_d_in_25_a),
    .io_d_in_25_valid_a(array_1_io_d_in_25_valid_a),
    .io_d_in_25_b(array_1_io_d_in_25_b),
    .io_d_in_25_valid_b(array_1_io_d_in_25_valid_b),
    .io_d_in_26_a(array_1_io_d_in_26_a),
    .io_d_in_26_valid_a(array_1_io_d_in_26_valid_a),
    .io_d_in_26_b(array_1_io_d_in_26_b),
    .io_d_in_26_valid_b(array_1_io_d_in_26_valid_b),
    .io_d_in_27_a(array_1_io_d_in_27_a),
    .io_d_in_27_valid_a(array_1_io_d_in_27_valid_a),
    .io_d_in_27_b(array_1_io_d_in_27_b),
    .io_d_in_27_valid_b(array_1_io_d_in_27_valid_b),
    .io_d_in_28_a(array_1_io_d_in_28_a),
    .io_d_in_28_valid_a(array_1_io_d_in_28_valid_a),
    .io_d_in_28_b(array_1_io_d_in_28_b),
    .io_d_in_28_valid_b(array_1_io_d_in_28_valid_b),
    .io_d_in_29_a(array_1_io_d_in_29_a),
    .io_d_in_29_valid_a(array_1_io_d_in_29_valid_a),
    .io_d_in_29_b(array_1_io_d_in_29_b),
    .io_d_in_29_valid_b(array_1_io_d_in_29_valid_b),
    .io_d_in_30_a(array_1_io_d_in_30_a),
    .io_d_in_30_valid_a(array_1_io_d_in_30_valid_a),
    .io_d_in_30_b(array_1_io_d_in_30_b),
    .io_d_in_30_valid_b(array_1_io_d_in_30_valid_b),
    .io_d_in_31_a(array_1_io_d_in_31_a),
    .io_d_in_31_valid_a(array_1_io_d_in_31_valid_a),
    .io_d_in_31_b(array_1_io_d_in_31_b),
    .io_d_in_31_valid_b(array_1_io_d_in_31_valid_b),
    .io_d_out_0_a(array_1_io_d_out_0_a),
    .io_d_out_0_valid_a(array_1_io_d_out_0_valid_a),
    .io_d_out_0_b(array_1_io_d_out_0_b),
    .io_d_out_0_valid_b(array_1_io_d_out_0_valid_b),
    .io_d_out_1_a(array_1_io_d_out_1_a),
    .io_d_out_1_valid_a(array_1_io_d_out_1_valid_a),
    .io_d_out_1_b(array_1_io_d_out_1_b),
    .io_d_out_1_valid_b(array_1_io_d_out_1_valid_b),
    .io_d_out_2_a(array_1_io_d_out_2_a),
    .io_d_out_2_valid_a(array_1_io_d_out_2_valid_a),
    .io_d_out_2_b(array_1_io_d_out_2_b),
    .io_d_out_2_valid_b(array_1_io_d_out_2_valid_b),
    .io_d_out_3_a(array_1_io_d_out_3_a),
    .io_d_out_3_valid_a(array_1_io_d_out_3_valid_a),
    .io_d_out_3_b(array_1_io_d_out_3_b),
    .io_d_out_3_valid_b(array_1_io_d_out_3_valid_b),
    .io_d_out_4_a(array_1_io_d_out_4_a),
    .io_d_out_4_valid_a(array_1_io_d_out_4_valid_a),
    .io_d_out_4_b(array_1_io_d_out_4_b),
    .io_d_out_4_valid_b(array_1_io_d_out_4_valid_b),
    .io_d_out_5_a(array_1_io_d_out_5_a),
    .io_d_out_5_valid_a(array_1_io_d_out_5_valid_a),
    .io_d_out_5_b(array_1_io_d_out_5_b),
    .io_d_out_5_valid_b(array_1_io_d_out_5_valid_b),
    .io_d_out_6_a(array_1_io_d_out_6_a),
    .io_d_out_6_valid_a(array_1_io_d_out_6_valid_a),
    .io_d_out_6_b(array_1_io_d_out_6_b),
    .io_d_out_6_valid_b(array_1_io_d_out_6_valid_b),
    .io_d_out_7_a(array_1_io_d_out_7_a),
    .io_d_out_7_valid_a(array_1_io_d_out_7_valid_a),
    .io_d_out_7_b(array_1_io_d_out_7_b),
    .io_d_out_7_valid_b(array_1_io_d_out_7_valid_b),
    .io_d_out_8_a(array_1_io_d_out_8_a),
    .io_d_out_8_valid_a(array_1_io_d_out_8_valid_a),
    .io_d_out_8_b(array_1_io_d_out_8_b),
    .io_d_out_8_valid_b(array_1_io_d_out_8_valid_b),
    .io_d_out_9_a(array_1_io_d_out_9_a),
    .io_d_out_9_valid_a(array_1_io_d_out_9_valid_a),
    .io_d_out_9_b(array_1_io_d_out_9_b),
    .io_d_out_9_valid_b(array_1_io_d_out_9_valid_b),
    .io_d_out_10_a(array_1_io_d_out_10_a),
    .io_d_out_10_valid_a(array_1_io_d_out_10_valid_a),
    .io_d_out_10_b(array_1_io_d_out_10_b),
    .io_d_out_10_valid_b(array_1_io_d_out_10_valid_b),
    .io_d_out_11_a(array_1_io_d_out_11_a),
    .io_d_out_11_valid_a(array_1_io_d_out_11_valid_a),
    .io_d_out_11_b(array_1_io_d_out_11_b),
    .io_d_out_11_valid_b(array_1_io_d_out_11_valid_b),
    .io_d_out_12_a(array_1_io_d_out_12_a),
    .io_d_out_12_valid_a(array_1_io_d_out_12_valid_a),
    .io_d_out_12_b(array_1_io_d_out_12_b),
    .io_d_out_12_valid_b(array_1_io_d_out_12_valid_b),
    .io_d_out_13_a(array_1_io_d_out_13_a),
    .io_d_out_13_valid_a(array_1_io_d_out_13_valid_a),
    .io_d_out_13_b(array_1_io_d_out_13_b),
    .io_d_out_13_valid_b(array_1_io_d_out_13_valid_b),
    .io_d_out_14_a(array_1_io_d_out_14_a),
    .io_d_out_14_valid_a(array_1_io_d_out_14_valid_a),
    .io_d_out_14_b(array_1_io_d_out_14_b),
    .io_d_out_14_valid_b(array_1_io_d_out_14_valid_b),
    .io_d_out_15_a(array_1_io_d_out_15_a),
    .io_d_out_15_valid_a(array_1_io_d_out_15_valid_a),
    .io_d_out_15_b(array_1_io_d_out_15_b),
    .io_d_out_15_valid_b(array_1_io_d_out_15_valid_b),
    .io_d_out_16_a(array_1_io_d_out_16_a),
    .io_d_out_16_valid_a(array_1_io_d_out_16_valid_a),
    .io_d_out_16_b(array_1_io_d_out_16_b),
    .io_d_out_16_valid_b(array_1_io_d_out_16_valid_b),
    .io_d_out_17_a(array_1_io_d_out_17_a),
    .io_d_out_17_valid_a(array_1_io_d_out_17_valid_a),
    .io_d_out_17_b(array_1_io_d_out_17_b),
    .io_d_out_17_valid_b(array_1_io_d_out_17_valid_b),
    .io_d_out_18_a(array_1_io_d_out_18_a),
    .io_d_out_18_valid_a(array_1_io_d_out_18_valid_a),
    .io_d_out_18_b(array_1_io_d_out_18_b),
    .io_d_out_18_valid_b(array_1_io_d_out_18_valid_b),
    .io_d_out_19_a(array_1_io_d_out_19_a),
    .io_d_out_19_valid_a(array_1_io_d_out_19_valid_a),
    .io_d_out_19_b(array_1_io_d_out_19_b),
    .io_d_out_19_valid_b(array_1_io_d_out_19_valid_b),
    .io_d_out_20_a(array_1_io_d_out_20_a),
    .io_d_out_20_valid_a(array_1_io_d_out_20_valid_a),
    .io_d_out_20_b(array_1_io_d_out_20_b),
    .io_d_out_20_valid_b(array_1_io_d_out_20_valid_b),
    .io_d_out_21_a(array_1_io_d_out_21_a),
    .io_d_out_21_valid_a(array_1_io_d_out_21_valid_a),
    .io_d_out_21_b(array_1_io_d_out_21_b),
    .io_d_out_21_valid_b(array_1_io_d_out_21_valid_b),
    .io_d_out_22_a(array_1_io_d_out_22_a),
    .io_d_out_22_valid_a(array_1_io_d_out_22_valid_a),
    .io_d_out_22_b(array_1_io_d_out_22_b),
    .io_d_out_22_valid_b(array_1_io_d_out_22_valid_b),
    .io_d_out_23_a(array_1_io_d_out_23_a),
    .io_d_out_23_valid_a(array_1_io_d_out_23_valid_a),
    .io_d_out_23_b(array_1_io_d_out_23_b),
    .io_d_out_23_valid_b(array_1_io_d_out_23_valid_b),
    .io_d_out_24_a(array_1_io_d_out_24_a),
    .io_d_out_24_valid_a(array_1_io_d_out_24_valid_a),
    .io_d_out_24_b(array_1_io_d_out_24_b),
    .io_d_out_24_valid_b(array_1_io_d_out_24_valid_b),
    .io_d_out_25_a(array_1_io_d_out_25_a),
    .io_d_out_25_valid_a(array_1_io_d_out_25_valid_a),
    .io_d_out_25_b(array_1_io_d_out_25_b),
    .io_d_out_25_valid_b(array_1_io_d_out_25_valid_b),
    .io_d_out_26_a(array_1_io_d_out_26_a),
    .io_d_out_26_valid_a(array_1_io_d_out_26_valid_a),
    .io_d_out_26_b(array_1_io_d_out_26_b),
    .io_d_out_26_valid_b(array_1_io_d_out_26_valid_b),
    .io_d_out_27_a(array_1_io_d_out_27_a),
    .io_d_out_27_valid_a(array_1_io_d_out_27_valid_a),
    .io_d_out_27_b(array_1_io_d_out_27_b),
    .io_d_out_27_valid_b(array_1_io_d_out_27_valid_b),
    .io_d_out_28_a(array_1_io_d_out_28_a),
    .io_d_out_28_valid_a(array_1_io_d_out_28_valid_a),
    .io_d_out_28_b(array_1_io_d_out_28_b),
    .io_d_out_28_valid_b(array_1_io_d_out_28_valid_b),
    .io_d_out_29_a(array_1_io_d_out_29_a),
    .io_d_out_29_valid_a(array_1_io_d_out_29_valid_a),
    .io_d_out_29_b(array_1_io_d_out_29_b),
    .io_d_out_29_valid_b(array_1_io_d_out_29_valid_b),
    .io_d_out_30_a(array_1_io_d_out_30_a),
    .io_d_out_30_valid_a(array_1_io_d_out_30_valid_a),
    .io_d_out_30_b(array_1_io_d_out_30_b),
    .io_d_out_30_valid_b(array_1_io_d_out_30_valid_b),
    .io_d_out_31_a(array_1_io_d_out_31_a),
    .io_d_out_31_valid_a(array_1_io_d_out_31_valid_a),
    .io_d_out_31_b(array_1_io_d_out_31_b),
    .io_d_out_31_valid_b(array_1_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_1_io_wr_en_mem1),
    .io_wr_en_mem2(array_1_io_wr_en_mem2),
    .io_wr_en_mem3(array_1_io_wr_en_mem3),
    .io_wr_en_mem4(array_1_io_wr_en_mem4),
    .io_wr_en_mem5(array_1_io_wr_en_mem5),
    .io_wr_en_mem6(array_1_io_wr_en_mem6),
    .io_wr_instr_mem1(array_1_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_1_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_1_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_1_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_1_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_1_io_wr_instr_mem6),
    .io_PC1_in(array_1_io_PC1_in),
    .io_PC6_out(array_1_io_PC6_out),
    .io_Addr_in(array_1_io_Addr_in),
    .io_Addr_out(array_1_io_Addr_out)
  );
  BuildingBlockNew array_2 ( // @[BP.scala 45:51]
    .clock(array_2_clock),
    .reset(array_2_reset),
    .io_d_in_0_a(array_2_io_d_in_0_a),
    .io_d_in_0_valid_a(array_2_io_d_in_0_valid_a),
    .io_d_in_0_b(array_2_io_d_in_0_b),
    .io_d_in_0_valid_b(array_2_io_d_in_0_valid_b),
    .io_d_in_1_a(array_2_io_d_in_1_a),
    .io_d_in_1_valid_a(array_2_io_d_in_1_valid_a),
    .io_d_in_1_b(array_2_io_d_in_1_b),
    .io_d_in_1_valid_b(array_2_io_d_in_1_valid_b),
    .io_d_in_2_a(array_2_io_d_in_2_a),
    .io_d_in_2_valid_a(array_2_io_d_in_2_valid_a),
    .io_d_in_2_b(array_2_io_d_in_2_b),
    .io_d_in_2_valid_b(array_2_io_d_in_2_valid_b),
    .io_d_in_3_a(array_2_io_d_in_3_a),
    .io_d_in_3_valid_a(array_2_io_d_in_3_valid_a),
    .io_d_in_3_b(array_2_io_d_in_3_b),
    .io_d_in_3_valid_b(array_2_io_d_in_3_valid_b),
    .io_d_in_4_a(array_2_io_d_in_4_a),
    .io_d_in_4_valid_a(array_2_io_d_in_4_valid_a),
    .io_d_in_4_b(array_2_io_d_in_4_b),
    .io_d_in_4_valid_b(array_2_io_d_in_4_valid_b),
    .io_d_in_5_a(array_2_io_d_in_5_a),
    .io_d_in_5_valid_a(array_2_io_d_in_5_valid_a),
    .io_d_in_5_b(array_2_io_d_in_5_b),
    .io_d_in_5_valid_b(array_2_io_d_in_5_valid_b),
    .io_d_in_6_a(array_2_io_d_in_6_a),
    .io_d_in_6_valid_a(array_2_io_d_in_6_valid_a),
    .io_d_in_6_b(array_2_io_d_in_6_b),
    .io_d_in_6_valid_b(array_2_io_d_in_6_valid_b),
    .io_d_in_7_a(array_2_io_d_in_7_a),
    .io_d_in_7_valid_a(array_2_io_d_in_7_valid_a),
    .io_d_in_7_b(array_2_io_d_in_7_b),
    .io_d_in_7_valid_b(array_2_io_d_in_7_valid_b),
    .io_d_in_8_a(array_2_io_d_in_8_a),
    .io_d_in_8_valid_a(array_2_io_d_in_8_valid_a),
    .io_d_in_8_b(array_2_io_d_in_8_b),
    .io_d_in_8_valid_b(array_2_io_d_in_8_valid_b),
    .io_d_in_9_a(array_2_io_d_in_9_a),
    .io_d_in_9_valid_a(array_2_io_d_in_9_valid_a),
    .io_d_in_9_b(array_2_io_d_in_9_b),
    .io_d_in_9_valid_b(array_2_io_d_in_9_valid_b),
    .io_d_in_10_a(array_2_io_d_in_10_a),
    .io_d_in_10_valid_a(array_2_io_d_in_10_valid_a),
    .io_d_in_10_b(array_2_io_d_in_10_b),
    .io_d_in_10_valid_b(array_2_io_d_in_10_valid_b),
    .io_d_in_11_a(array_2_io_d_in_11_a),
    .io_d_in_11_valid_a(array_2_io_d_in_11_valid_a),
    .io_d_in_11_b(array_2_io_d_in_11_b),
    .io_d_in_11_valid_b(array_2_io_d_in_11_valid_b),
    .io_d_in_12_a(array_2_io_d_in_12_a),
    .io_d_in_12_valid_a(array_2_io_d_in_12_valid_a),
    .io_d_in_12_b(array_2_io_d_in_12_b),
    .io_d_in_12_valid_b(array_2_io_d_in_12_valid_b),
    .io_d_in_13_a(array_2_io_d_in_13_a),
    .io_d_in_13_valid_a(array_2_io_d_in_13_valid_a),
    .io_d_in_13_b(array_2_io_d_in_13_b),
    .io_d_in_13_valid_b(array_2_io_d_in_13_valid_b),
    .io_d_in_14_a(array_2_io_d_in_14_a),
    .io_d_in_14_valid_a(array_2_io_d_in_14_valid_a),
    .io_d_in_14_b(array_2_io_d_in_14_b),
    .io_d_in_14_valid_b(array_2_io_d_in_14_valid_b),
    .io_d_in_15_a(array_2_io_d_in_15_a),
    .io_d_in_15_valid_a(array_2_io_d_in_15_valid_a),
    .io_d_in_15_b(array_2_io_d_in_15_b),
    .io_d_in_15_valid_b(array_2_io_d_in_15_valid_b),
    .io_d_in_16_a(array_2_io_d_in_16_a),
    .io_d_in_16_valid_a(array_2_io_d_in_16_valid_a),
    .io_d_in_16_b(array_2_io_d_in_16_b),
    .io_d_in_16_valid_b(array_2_io_d_in_16_valid_b),
    .io_d_in_17_a(array_2_io_d_in_17_a),
    .io_d_in_17_valid_a(array_2_io_d_in_17_valid_a),
    .io_d_in_17_b(array_2_io_d_in_17_b),
    .io_d_in_17_valid_b(array_2_io_d_in_17_valid_b),
    .io_d_in_18_a(array_2_io_d_in_18_a),
    .io_d_in_18_valid_a(array_2_io_d_in_18_valid_a),
    .io_d_in_18_b(array_2_io_d_in_18_b),
    .io_d_in_18_valid_b(array_2_io_d_in_18_valid_b),
    .io_d_in_19_a(array_2_io_d_in_19_a),
    .io_d_in_19_valid_a(array_2_io_d_in_19_valid_a),
    .io_d_in_19_b(array_2_io_d_in_19_b),
    .io_d_in_19_valid_b(array_2_io_d_in_19_valid_b),
    .io_d_in_20_a(array_2_io_d_in_20_a),
    .io_d_in_20_valid_a(array_2_io_d_in_20_valid_a),
    .io_d_in_20_b(array_2_io_d_in_20_b),
    .io_d_in_20_valid_b(array_2_io_d_in_20_valid_b),
    .io_d_in_21_a(array_2_io_d_in_21_a),
    .io_d_in_21_valid_a(array_2_io_d_in_21_valid_a),
    .io_d_in_21_b(array_2_io_d_in_21_b),
    .io_d_in_21_valid_b(array_2_io_d_in_21_valid_b),
    .io_d_in_22_a(array_2_io_d_in_22_a),
    .io_d_in_22_valid_a(array_2_io_d_in_22_valid_a),
    .io_d_in_22_b(array_2_io_d_in_22_b),
    .io_d_in_22_valid_b(array_2_io_d_in_22_valid_b),
    .io_d_in_23_a(array_2_io_d_in_23_a),
    .io_d_in_23_valid_a(array_2_io_d_in_23_valid_a),
    .io_d_in_23_b(array_2_io_d_in_23_b),
    .io_d_in_23_valid_b(array_2_io_d_in_23_valid_b),
    .io_d_in_24_a(array_2_io_d_in_24_a),
    .io_d_in_24_valid_a(array_2_io_d_in_24_valid_a),
    .io_d_in_24_b(array_2_io_d_in_24_b),
    .io_d_in_24_valid_b(array_2_io_d_in_24_valid_b),
    .io_d_in_25_a(array_2_io_d_in_25_a),
    .io_d_in_25_valid_a(array_2_io_d_in_25_valid_a),
    .io_d_in_25_b(array_2_io_d_in_25_b),
    .io_d_in_25_valid_b(array_2_io_d_in_25_valid_b),
    .io_d_in_26_a(array_2_io_d_in_26_a),
    .io_d_in_26_valid_a(array_2_io_d_in_26_valid_a),
    .io_d_in_26_b(array_2_io_d_in_26_b),
    .io_d_in_26_valid_b(array_2_io_d_in_26_valid_b),
    .io_d_in_27_a(array_2_io_d_in_27_a),
    .io_d_in_27_valid_a(array_2_io_d_in_27_valid_a),
    .io_d_in_27_b(array_2_io_d_in_27_b),
    .io_d_in_27_valid_b(array_2_io_d_in_27_valid_b),
    .io_d_in_28_a(array_2_io_d_in_28_a),
    .io_d_in_28_valid_a(array_2_io_d_in_28_valid_a),
    .io_d_in_28_b(array_2_io_d_in_28_b),
    .io_d_in_28_valid_b(array_2_io_d_in_28_valid_b),
    .io_d_in_29_a(array_2_io_d_in_29_a),
    .io_d_in_29_valid_a(array_2_io_d_in_29_valid_a),
    .io_d_in_29_b(array_2_io_d_in_29_b),
    .io_d_in_29_valid_b(array_2_io_d_in_29_valid_b),
    .io_d_in_30_a(array_2_io_d_in_30_a),
    .io_d_in_30_valid_a(array_2_io_d_in_30_valid_a),
    .io_d_in_30_b(array_2_io_d_in_30_b),
    .io_d_in_30_valid_b(array_2_io_d_in_30_valid_b),
    .io_d_in_31_a(array_2_io_d_in_31_a),
    .io_d_in_31_valid_a(array_2_io_d_in_31_valid_a),
    .io_d_in_31_b(array_2_io_d_in_31_b),
    .io_d_in_31_valid_b(array_2_io_d_in_31_valid_b),
    .io_d_out_0_a(array_2_io_d_out_0_a),
    .io_d_out_0_valid_a(array_2_io_d_out_0_valid_a),
    .io_d_out_0_b(array_2_io_d_out_0_b),
    .io_d_out_0_valid_b(array_2_io_d_out_0_valid_b),
    .io_d_out_1_a(array_2_io_d_out_1_a),
    .io_d_out_1_valid_a(array_2_io_d_out_1_valid_a),
    .io_d_out_1_b(array_2_io_d_out_1_b),
    .io_d_out_1_valid_b(array_2_io_d_out_1_valid_b),
    .io_d_out_2_a(array_2_io_d_out_2_a),
    .io_d_out_2_valid_a(array_2_io_d_out_2_valid_a),
    .io_d_out_2_b(array_2_io_d_out_2_b),
    .io_d_out_2_valid_b(array_2_io_d_out_2_valid_b),
    .io_d_out_3_a(array_2_io_d_out_3_a),
    .io_d_out_3_valid_a(array_2_io_d_out_3_valid_a),
    .io_d_out_3_b(array_2_io_d_out_3_b),
    .io_d_out_3_valid_b(array_2_io_d_out_3_valid_b),
    .io_d_out_4_a(array_2_io_d_out_4_a),
    .io_d_out_4_valid_a(array_2_io_d_out_4_valid_a),
    .io_d_out_4_b(array_2_io_d_out_4_b),
    .io_d_out_4_valid_b(array_2_io_d_out_4_valid_b),
    .io_d_out_5_a(array_2_io_d_out_5_a),
    .io_d_out_5_valid_a(array_2_io_d_out_5_valid_a),
    .io_d_out_5_b(array_2_io_d_out_5_b),
    .io_d_out_5_valid_b(array_2_io_d_out_5_valid_b),
    .io_d_out_6_a(array_2_io_d_out_6_a),
    .io_d_out_6_valid_a(array_2_io_d_out_6_valid_a),
    .io_d_out_6_b(array_2_io_d_out_6_b),
    .io_d_out_6_valid_b(array_2_io_d_out_6_valid_b),
    .io_d_out_7_a(array_2_io_d_out_7_a),
    .io_d_out_7_valid_a(array_2_io_d_out_7_valid_a),
    .io_d_out_7_b(array_2_io_d_out_7_b),
    .io_d_out_7_valid_b(array_2_io_d_out_7_valid_b),
    .io_d_out_8_a(array_2_io_d_out_8_a),
    .io_d_out_8_valid_a(array_2_io_d_out_8_valid_a),
    .io_d_out_8_b(array_2_io_d_out_8_b),
    .io_d_out_8_valid_b(array_2_io_d_out_8_valid_b),
    .io_d_out_9_a(array_2_io_d_out_9_a),
    .io_d_out_9_valid_a(array_2_io_d_out_9_valid_a),
    .io_d_out_9_b(array_2_io_d_out_9_b),
    .io_d_out_9_valid_b(array_2_io_d_out_9_valid_b),
    .io_d_out_10_a(array_2_io_d_out_10_a),
    .io_d_out_10_valid_a(array_2_io_d_out_10_valid_a),
    .io_d_out_10_b(array_2_io_d_out_10_b),
    .io_d_out_10_valid_b(array_2_io_d_out_10_valid_b),
    .io_d_out_11_a(array_2_io_d_out_11_a),
    .io_d_out_11_valid_a(array_2_io_d_out_11_valid_a),
    .io_d_out_11_b(array_2_io_d_out_11_b),
    .io_d_out_11_valid_b(array_2_io_d_out_11_valid_b),
    .io_d_out_12_a(array_2_io_d_out_12_a),
    .io_d_out_12_valid_a(array_2_io_d_out_12_valid_a),
    .io_d_out_12_b(array_2_io_d_out_12_b),
    .io_d_out_12_valid_b(array_2_io_d_out_12_valid_b),
    .io_d_out_13_a(array_2_io_d_out_13_a),
    .io_d_out_13_valid_a(array_2_io_d_out_13_valid_a),
    .io_d_out_13_b(array_2_io_d_out_13_b),
    .io_d_out_13_valid_b(array_2_io_d_out_13_valid_b),
    .io_d_out_14_a(array_2_io_d_out_14_a),
    .io_d_out_14_valid_a(array_2_io_d_out_14_valid_a),
    .io_d_out_14_b(array_2_io_d_out_14_b),
    .io_d_out_14_valid_b(array_2_io_d_out_14_valid_b),
    .io_d_out_15_a(array_2_io_d_out_15_a),
    .io_d_out_15_valid_a(array_2_io_d_out_15_valid_a),
    .io_d_out_15_b(array_2_io_d_out_15_b),
    .io_d_out_15_valid_b(array_2_io_d_out_15_valid_b),
    .io_d_out_16_a(array_2_io_d_out_16_a),
    .io_d_out_16_valid_a(array_2_io_d_out_16_valid_a),
    .io_d_out_16_b(array_2_io_d_out_16_b),
    .io_d_out_16_valid_b(array_2_io_d_out_16_valid_b),
    .io_d_out_17_a(array_2_io_d_out_17_a),
    .io_d_out_17_valid_a(array_2_io_d_out_17_valid_a),
    .io_d_out_17_b(array_2_io_d_out_17_b),
    .io_d_out_17_valid_b(array_2_io_d_out_17_valid_b),
    .io_d_out_18_a(array_2_io_d_out_18_a),
    .io_d_out_18_valid_a(array_2_io_d_out_18_valid_a),
    .io_d_out_18_b(array_2_io_d_out_18_b),
    .io_d_out_18_valid_b(array_2_io_d_out_18_valid_b),
    .io_d_out_19_a(array_2_io_d_out_19_a),
    .io_d_out_19_valid_a(array_2_io_d_out_19_valid_a),
    .io_d_out_19_b(array_2_io_d_out_19_b),
    .io_d_out_19_valid_b(array_2_io_d_out_19_valid_b),
    .io_d_out_20_a(array_2_io_d_out_20_a),
    .io_d_out_20_valid_a(array_2_io_d_out_20_valid_a),
    .io_d_out_20_b(array_2_io_d_out_20_b),
    .io_d_out_20_valid_b(array_2_io_d_out_20_valid_b),
    .io_d_out_21_a(array_2_io_d_out_21_a),
    .io_d_out_21_valid_a(array_2_io_d_out_21_valid_a),
    .io_d_out_21_b(array_2_io_d_out_21_b),
    .io_d_out_21_valid_b(array_2_io_d_out_21_valid_b),
    .io_d_out_22_a(array_2_io_d_out_22_a),
    .io_d_out_22_valid_a(array_2_io_d_out_22_valid_a),
    .io_d_out_22_b(array_2_io_d_out_22_b),
    .io_d_out_22_valid_b(array_2_io_d_out_22_valid_b),
    .io_d_out_23_a(array_2_io_d_out_23_a),
    .io_d_out_23_valid_a(array_2_io_d_out_23_valid_a),
    .io_d_out_23_b(array_2_io_d_out_23_b),
    .io_d_out_23_valid_b(array_2_io_d_out_23_valid_b),
    .io_d_out_24_a(array_2_io_d_out_24_a),
    .io_d_out_24_valid_a(array_2_io_d_out_24_valid_a),
    .io_d_out_24_b(array_2_io_d_out_24_b),
    .io_d_out_24_valid_b(array_2_io_d_out_24_valid_b),
    .io_d_out_25_a(array_2_io_d_out_25_a),
    .io_d_out_25_valid_a(array_2_io_d_out_25_valid_a),
    .io_d_out_25_b(array_2_io_d_out_25_b),
    .io_d_out_25_valid_b(array_2_io_d_out_25_valid_b),
    .io_d_out_26_a(array_2_io_d_out_26_a),
    .io_d_out_26_valid_a(array_2_io_d_out_26_valid_a),
    .io_d_out_26_b(array_2_io_d_out_26_b),
    .io_d_out_26_valid_b(array_2_io_d_out_26_valid_b),
    .io_d_out_27_a(array_2_io_d_out_27_a),
    .io_d_out_27_valid_a(array_2_io_d_out_27_valid_a),
    .io_d_out_27_b(array_2_io_d_out_27_b),
    .io_d_out_27_valid_b(array_2_io_d_out_27_valid_b),
    .io_d_out_28_a(array_2_io_d_out_28_a),
    .io_d_out_28_valid_a(array_2_io_d_out_28_valid_a),
    .io_d_out_28_b(array_2_io_d_out_28_b),
    .io_d_out_28_valid_b(array_2_io_d_out_28_valid_b),
    .io_d_out_29_a(array_2_io_d_out_29_a),
    .io_d_out_29_valid_a(array_2_io_d_out_29_valid_a),
    .io_d_out_29_b(array_2_io_d_out_29_b),
    .io_d_out_29_valid_b(array_2_io_d_out_29_valid_b),
    .io_d_out_30_a(array_2_io_d_out_30_a),
    .io_d_out_30_valid_a(array_2_io_d_out_30_valid_a),
    .io_d_out_30_b(array_2_io_d_out_30_b),
    .io_d_out_30_valid_b(array_2_io_d_out_30_valid_b),
    .io_d_out_31_a(array_2_io_d_out_31_a),
    .io_d_out_31_valid_a(array_2_io_d_out_31_valid_a),
    .io_d_out_31_b(array_2_io_d_out_31_b),
    .io_d_out_31_valid_b(array_2_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_2_io_wr_en_mem1),
    .io_wr_en_mem2(array_2_io_wr_en_mem2),
    .io_wr_en_mem3(array_2_io_wr_en_mem3),
    .io_wr_en_mem4(array_2_io_wr_en_mem4),
    .io_wr_en_mem5(array_2_io_wr_en_mem5),
    .io_wr_en_mem6(array_2_io_wr_en_mem6),
    .io_wr_instr_mem1(array_2_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_2_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_2_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_2_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_2_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_2_io_wr_instr_mem6),
    .io_PC1_in(array_2_io_PC1_in),
    .io_PC6_out(array_2_io_PC6_out),
    .io_Addr_in(array_2_io_Addr_in),
    .io_Addr_out(array_2_io_Addr_out)
  );
  BuildingBlockNew array_3 ( // @[BP.scala 45:51]
    .clock(array_3_clock),
    .reset(array_3_reset),
    .io_d_in_0_a(array_3_io_d_in_0_a),
    .io_d_in_0_valid_a(array_3_io_d_in_0_valid_a),
    .io_d_in_0_b(array_3_io_d_in_0_b),
    .io_d_in_0_valid_b(array_3_io_d_in_0_valid_b),
    .io_d_in_1_a(array_3_io_d_in_1_a),
    .io_d_in_1_valid_a(array_3_io_d_in_1_valid_a),
    .io_d_in_1_b(array_3_io_d_in_1_b),
    .io_d_in_1_valid_b(array_3_io_d_in_1_valid_b),
    .io_d_in_2_a(array_3_io_d_in_2_a),
    .io_d_in_2_valid_a(array_3_io_d_in_2_valid_a),
    .io_d_in_2_b(array_3_io_d_in_2_b),
    .io_d_in_2_valid_b(array_3_io_d_in_2_valid_b),
    .io_d_in_3_a(array_3_io_d_in_3_a),
    .io_d_in_3_valid_a(array_3_io_d_in_3_valid_a),
    .io_d_in_3_b(array_3_io_d_in_3_b),
    .io_d_in_3_valid_b(array_3_io_d_in_3_valid_b),
    .io_d_in_4_a(array_3_io_d_in_4_a),
    .io_d_in_4_valid_a(array_3_io_d_in_4_valid_a),
    .io_d_in_4_b(array_3_io_d_in_4_b),
    .io_d_in_4_valid_b(array_3_io_d_in_4_valid_b),
    .io_d_in_5_a(array_3_io_d_in_5_a),
    .io_d_in_5_valid_a(array_3_io_d_in_5_valid_a),
    .io_d_in_5_b(array_3_io_d_in_5_b),
    .io_d_in_5_valid_b(array_3_io_d_in_5_valid_b),
    .io_d_in_6_a(array_3_io_d_in_6_a),
    .io_d_in_6_valid_a(array_3_io_d_in_6_valid_a),
    .io_d_in_6_b(array_3_io_d_in_6_b),
    .io_d_in_6_valid_b(array_3_io_d_in_6_valid_b),
    .io_d_in_7_a(array_3_io_d_in_7_a),
    .io_d_in_7_valid_a(array_3_io_d_in_7_valid_a),
    .io_d_in_7_b(array_3_io_d_in_7_b),
    .io_d_in_7_valid_b(array_3_io_d_in_7_valid_b),
    .io_d_in_8_a(array_3_io_d_in_8_a),
    .io_d_in_8_valid_a(array_3_io_d_in_8_valid_a),
    .io_d_in_8_b(array_3_io_d_in_8_b),
    .io_d_in_8_valid_b(array_3_io_d_in_8_valid_b),
    .io_d_in_9_a(array_3_io_d_in_9_a),
    .io_d_in_9_valid_a(array_3_io_d_in_9_valid_a),
    .io_d_in_9_b(array_3_io_d_in_9_b),
    .io_d_in_9_valid_b(array_3_io_d_in_9_valid_b),
    .io_d_in_10_a(array_3_io_d_in_10_a),
    .io_d_in_10_valid_a(array_3_io_d_in_10_valid_a),
    .io_d_in_10_b(array_3_io_d_in_10_b),
    .io_d_in_10_valid_b(array_3_io_d_in_10_valid_b),
    .io_d_in_11_a(array_3_io_d_in_11_a),
    .io_d_in_11_valid_a(array_3_io_d_in_11_valid_a),
    .io_d_in_11_b(array_3_io_d_in_11_b),
    .io_d_in_11_valid_b(array_3_io_d_in_11_valid_b),
    .io_d_in_12_a(array_3_io_d_in_12_a),
    .io_d_in_12_valid_a(array_3_io_d_in_12_valid_a),
    .io_d_in_12_b(array_3_io_d_in_12_b),
    .io_d_in_12_valid_b(array_3_io_d_in_12_valid_b),
    .io_d_in_13_a(array_3_io_d_in_13_a),
    .io_d_in_13_valid_a(array_3_io_d_in_13_valid_a),
    .io_d_in_13_b(array_3_io_d_in_13_b),
    .io_d_in_13_valid_b(array_3_io_d_in_13_valid_b),
    .io_d_in_14_a(array_3_io_d_in_14_a),
    .io_d_in_14_valid_a(array_3_io_d_in_14_valid_a),
    .io_d_in_14_b(array_3_io_d_in_14_b),
    .io_d_in_14_valid_b(array_3_io_d_in_14_valid_b),
    .io_d_in_15_a(array_3_io_d_in_15_a),
    .io_d_in_15_valid_a(array_3_io_d_in_15_valid_a),
    .io_d_in_15_b(array_3_io_d_in_15_b),
    .io_d_in_15_valid_b(array_3_io_d_in_15_valid_b),
    .io_d_in_16_a(array_3_io_d_in_16_a),
    .io_d_in_16_valid_a(array_3_io_d_in_16_valid_a),
    .io_d_in_16_b(array_3_io_d_in_16_b),
    .io_d_in_16_valid_b(array_3_io_d_in_16_valid_b),
    .io_d_in_17_a(array_3_io_d_in_17_a),
    .io_d_in_17_valid_a(array_3_io_d_in_17_valid_a),
    .io_d_in_17_b(array_3_io_d_in_17_b),
    .io_d_in_17_valid_b(array_3_io_d_in_17_valid_b),
    .io_d_in_18_a(array_3_io_d_in_18_a),
    .io_d_in_18_valid_a(array_3_io_d_in_18_valid_a),
    .io_d_in_18_b(array_3_io_d_in_18_b),
    .io_d_in_18_valid_b(array_3_io_d_in_18_valid_b),
    .io_d_in_19_a(array_3_io_d_in_19_a),
    .io_d_in_19_valid_a(array_3_io_d_in_19_valid_a),
    .io_d_in_19_b(array_3_io_d_in_19_b),
    .io_d_in_19_valid_b(array_3_io_d_in_19_valid_b),
    .io_d_in_20_a(array_3_io_d_in_20_a),
    .io_d_in_20_valid_a(array_3_io_d_in_20_valid_a),
    .io_d_in_20_b(array_3_io_d_in_20_b),
    .io_d_in_20_valid_b(array_3_io_d_in_20_valid_b),
    .io_d_in_21_a(array_3_io_d_in_21_a),
    .io_d_in_21_valid_a(array_3_io_d_in_21_valid_a),
    .io_d_in_21_b(array_3_io_d_in_21_b),
    .io_d_in_21_valid_b(array_3_io_d_in_21_valid_b),
    .io_d_in_22_a(array_3_io_d_in_22_a),
    .io_d_in_22_valid_a(array_3_io_d_in_22_valid_a),
    .io_d_in_22_b(array_3_io_d_in_22_b),
    .io_d_in_22_valid_b(array_3_io_d_in_22_valid_b),
    .io_d_in_23_a(array_3_io_d_in_23_a),
    .io_d_in_23_valid_a(array_3_io_d_in_23_valid_a),
    .io_d_in_23_b(array_3_io_d_in_23_b),
    .io_d_in_23_valid_b(array_3_io_d_in_23_valid_b),
    .io_d_in_24_a(array_3_io_d_in_24_a),
    .io_d_in_24_valid_a(array_3_io_d_in_24_valid_a),
    .io_d_in_24_b(array_3_io_d_in_24_b),
    .io_d_in_24_valid_b(array_3_io_d_in_24_valid_b),
    .io_d_in_25_a(array_3_io_d_in_25_a),
    .io_d_in_25_valid_a(array_3_io_d_in_25_valid_a),
    .io_d_in_25_b(array_3_io_d_in_25_b),
    .io_d_in_25_valid_b(array_3_io_d_in_25_valid_b),
    .io_d_in_26_a(array_3_io_d_in_26_a),
    .io_d_in_26_valid_a(array_3_io_d_in_26_valid_a),
    .io_d_in_26_b(array_3_io_d_in_26_b),
    .io_d_in_26_valid_b(array_3_io_d_in_26_valid_b),
    .io_d_in_27_a(array_3_io_d_in_27_a),
    .io_d_in_27_valid_a(array_3_io_d_in_27_valid_a),
    .io_d_in_27_b(array_3_io_d_in_27_b),
    .io_d_in_27_valid_b(array_3_io_d_in_27_valid_b),
    .io_d_in_28_a(array_3_io_d_in_28_a),
    .io_d_in_28_valid_a(array_3_io_d_in_28_valid_a),
    .io_d_in_28_b(array_3_io_d_in_28_b),
    .io_d_in_28_valid_b(array_3_io_d_in_28_valid_b),
    .io_d_in_29_a(array_3_io_d_in_29_a),
    .io_d_in_29_valid_a(array_3_io_d_in_29_valid_a),
    .io_d_in_29_b(array_3_io_d_in_29_b),
    .io_d_in_29_valid_b(array_3_io_d_in_29_valid_b),
    .io_d_in_30_a(array_3_io_d_in_30_a),
    .io_d_in_30_valid_a(array_3_io_d_in_30_valid_a),
    .io_d_in_30_b(array_3_io_d_in_30_b),
    .io_d_in_30_valid_b(array_3_io_d_in_30_valid_b),
    .io_d_in_31_a(array_3_io_d_in_31_a),
    .io_d_in_31_valid_a(array_3_io_d_in_31_valid_a),
    .io_d_in_31_b(array_3_io_d_in_31_b),
    .io_d_in_31_valid_b(array_3_io_d_in_31_valid_b),
    .io_d_out_0_a(array_3_io_d_out_0_a),
    .io_d_out_0_valid_a(array_3_io_d_out_0_valid_a),
    .io_d_out_0_b(array_3_io_d_out_0_b),
    .io_d_out_0_valid_b(array_3_io_d_out_0_valid_b),
    .io_d_out_1_a(array_3_io_d_out_1_a),
    .io_d_out_1_valid_a(array_3_io_d_out_1_valid_a),
    .io_d_out_1_b(array_3_io_d_out_1_b),
    .io_d_out_1_valid_b(array_3_io_d_out_1_valid_b),
    .io_d_out_2_a(array_3_io_d_out_2_a),
    .io_d_out_2_valid_a(array_3_io_d_out_2_valid_a),
    .io_d_out_2_b(array_3_io_d_out_2_b),
    .io_d_out_2_valid_b(array_3_io_d_out_2_valid_b),
    .io_d_out_3_a(array_3_io_d_out_3_a),
    .io_d_out_3_valid_a(array_3_io_d_out_3_valid_a),
    .io_d_out_3_b(array_3_io_d_out_3_b),
    .io_d_out_3_valid_b(array_3_io_d_out_3_valid_b),
    .io_d_out_4_a(array_3_io_d_out_4_a),
    .io_d_out_4_valid_a(array_3_io_d_out_4_valid_a),
    .io_d_out_4_b(array_3_io_d_out_4_b),
    .io_d_out_4_valid_b(array_3_io_d_out_4_valid_b),
    .io_d_out_5_a(array_3_io_d_out_5_a),
    .io_d_out_5_valid_a(array_3_io_d_out_5_valid_a),
    .io_d_out_5_b(array_3_io_d_out_5_b),
    .io_d_out_5_valid_b(array_3_io_d_out_5_valid_b),
    .io_d_out_6_a(array_3_io_d_out_6_a),
    .io_d_out_6_valid_a(array_3_io_d_out_6_valid_a),
    .io_d_out_6_b(array_3_io_d_out_6_b),
    .io_d_out_6_valid_b(array_3_io_d_out_6_valid_b),
    .io_d_out_7_a(array_3_io_d_out_7_a),
    .io_d_out_7_valid_a(array_3_io_d_out_7_valid_a),
    .io_d_out_7_b(array_3_io_d_out_7_b),
    .io_d_out_7_valid_b(array_3_io_d_out_7_valid_b),
    .io_d_out_8_a(array_3_io_d_out_8_a),
    .io_d_out_8_valid_a(array_3_io_d_out_8_valid_a),
    .io_d_out_8_b(array_3_io_d_out_8_b),
    .io_d_out_8_valid_b(array_3_io_d_out_8_valid_b),
    .io_d_out_9_a(array_3_io_d_out_9_a),
    .io_d_out_9_valid_a(array_3_io_d_out_9_valid_a),
    .io_d_out_9_b(array_3_io_d_out_9_b),
    .io_d_out_9_valid_b(array_3_io_d_out_9_valid_b),
    .io_d_out_10_a(array_3_io_d_out_10_a),
    .io_d_out_10_valid_a(array_3_io_d_out_10_valid_a),
    .io_d_out_10_b(array_3_io_d_out_10_b),
    .io_d_out_10_valid_b(array_3_io_d_out_10_valid_b),
    .io_d_out_11_a(array_3_io_d_out_11_a),
    .io_d_out_11_valid_a(array_3_io_d_out_11_valid_a),
    .io_d_out_11_b(array_3_io_d_out_11_b),
    .io_d_out_11_valid_b(array_3_io_d_out_11_valid_b),
    .io_d_out_12_a(array_3_io_d_out_12_a),
    .io_d_out_12_valid_a(array_3_io_d_out_12_valid_a),
    .io_d_out_12_b(array_3_io_d_out_12_b),
    .io_d_out_12_valid_b(array_3_io_d_out_12_valid_b),
    .io_d_out_13_a(array_3_io_d_out_13_a),
    .io_d_out_13_valid_a(array_3_io_d_out_13_valid_a),
    .io_d_out_13_b(array_3_io_d_out_13_b),
    .io_d_out_13_valid_b(array_3_io_d_out_13_valid_b),
    .io_d_out_14_a(array_3_io_d_out_14_a),
    .io_d_out_14_valid_a(array_3_io_d_out_14_valid_a),
    .io_d_out_14_b(array_3_io_d_out_14_b),
    .io_d_out_14_valid_b(array_3_io_d_out_14_valid_b),
    .io_d_out_15_a(array_3_io_d_out_15_a),
    .io_d_out_15_valid_a(array_3_io_d_out_15_valid_a),
    .io_d_out_15_b(array_3_io_d_out_15_b),
    .io_d_out_15_valid_b(array_3_io_d_out_15_valid_b),
    .io_d_out_16_a(array_3_io_d_out_16_a),
    .io_d_out_16_valid_a(array_3_io_d_out_16_valid_a),
    .io_d_out_16_b(array_3_io_d_out_16_b),
    .io_d_out_16_valid_b(array_3_io_d_out_16_valid_b),
    .io_d_out_17_a(array_3_io_d_out_17_a),
    .io_d_out_17_valid_a(array_3_io_d_out_17_valid_a),
    .io_d_out_17_b(array_3_io_d_out_17_b),
    .io_d_out_17_valid_b(array_3_io_d_out_17_valid_b),
    .io_d_out_18_a(array_3_io_d_out_18_a),
    .io_d_out_18_valid_a(array_3_io_d_out_18_valid_a),
    .io_d_out_18_b(array_3_io_d_out_18_b),
    .io_d_out_18_valid_b(array_3_io_d_out_18_valid_b),
    .io_d_out_19_a(array_3_io_d_out_19_a),
    .io_d_out_19_valid_a(array_3_io_d_out_19_valid_a),
    .io_d_out_19_b(array_3_io_d_out_19_b),
    .io_d_out_19_valid_b(array_3_io_d_out_19_valid_b),
    .io_d_out_20_a(array_3_io_d_out_20_a),
    .io_d_out_20_valid_a(array_3_io_d_out_20_valid_a),
    .io_d_out_20_b(array_3_io_d_out_20_b),
    .io_d_out_20_valid_b(array_3_io_d_out_20_valid_b),
    .io_d_out_21_a(array_3_io_d_out_21_a),
    .io_d_out_21_valid_a(array_3_io_d_out_21_valid_a),
    .io_d_out_21_b(array_3_io_d_out_21_b),
    .io_d_out_21_valid_b(array_3_io_d_out_21_valid_b),
    .io_d_out_22_a(array_3_io_d_out_22_a),
    .io_d_out_22_valid_a(array_3_io_d_out_22_valid_a),
    .io_d_out_22_b(array_3_io_d_out_22_b),
    .io_d_out_22_valid_b(array_3_io_d_out_22_valid_b),
    .io_d_out_23_a(array_3_io_d_out_23_a),
    .io_d_out_23_valid_a(array_3_io_d_out_23_valid_a),
    .io_d_out_23_b(array_3_io_d_out_23_b),
    .io_d_out_23_valid_b(array_3_io_d_out_23_valid_b),
    .io_d_out_24_a(array_3_io_d_out_24_a),
    .io_d_out_24_valid_a(array_3_io_d_out_24_valid_a),
    .io_d_out_24_b(array_3_io_d_out_24_b),
    .io_d_out_24_valid_b(array_3_io_d_out_24_valid_b),
    .io_d_out_25_a(array_3_io_d_out_25_a),
    .io_d_out_25_valid_a(array_3_io_d_out_25_valid_a),
    .io_d_out_25_b(array_3_io_d_out_25_b),
    .io_d_out_25_valid_b(array_3_io_d_out_25_valid_b),
    .io_d_out_26_a(array_3_io_d_out_26_a),
    .io_d_out_26_valid_a(array_3_io_d_out_26_valid_a),
    .io_d_out_26_b(array_3_io_d_out_26_b),
    .io_d_out_26_valid_b(array_3_io_d_out_26_valid_b),
    .io_d_out_27_a(array_3_io_d_out_27_a),
    .io_d_out_27_valid_a(array_3_io_d_out_27_valid_a),
    .io_d_out_27_b(array_3_io_d_out_27_b),
    .io_d_out_27_valid_b(array_3_io_d_out_27_valid_b),
    .io_d_out_28_a(array_3_io_d_out_28_a),
    .io_d_out_28_valid_a(array_3_io_d_out_28_valid_a),
    .io_d_out_28_b(array_3_io_d_out_28_b),
    .io_d_out_28_valid_b(array_3_io_d_out_28_valid_b),
    .io_d_out_29_a(array_3_io_d_out_29_a),
    .io_d_out_29_valid_a(array_3_io_d_out_29_valid_a),
    .io_d_out_29_b(array_3_io_d_out_29_b),
    .io_d_out_29_valid_b(array_3_io_d_out_29_valid_b),
    .io_d_out_30_a(array_3_io_d_out_30_a),
    .io_d_out_30_valid_a(array_3_io_d_out_30_valid_a),
    .io_d_out_30_b(array_3_io_d_out_30_b),
    .io_d_out_30_valid_b(array_3_io_d_out_30_valid_b),
    .io_d_out_31_a(array_3_io_d_out_31_a),
    .io_d_out_31_valid_a(array_3_io_d_out_31_valid_a),
    .io_d_out_31_b(array_3_io_d_out_31_b),
    .io_d_out_31_valid_b(array_3_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_3_io_wr_en_mem1),
    .io_wr_en_mem2(array_3_io_wr_en_mem2),
    .io_wr_en_mem3(array_3_io_wr_en_mem3),
    .io_wr_en_mem4(array_3_io_wr_en_mem4),
    .io_wr_en_mem5(array_3_io_wr_en_mem5),
    .io_wr_en_mem6(array_3_io_wr_en_mem6),
    .io_wr_instr_mem1(array_3_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_3_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_3_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_3_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_3_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_3_io_wr_instr_mem6),
    .io_PC1_in(array_3_io_PC1_in),
    .io_PC6_out(array_3_io_PC6_out),
    .io_Addr_in(array_3_io_Addr_in),
    .io_Addr_out(array_3_io_Addr_out)
  );
  BuildingBlockNew array_4 ( // @[BP.scala 45:51]
    .clock(array_4_clock),
    .reset(array_4_reset),
    .io_d_in_0_a(array_4_io_d_in_0_a),
    .io_d_in_0_valid_a(array_4_io_d_in_0_valid_a),
    .io_d_in_0_b(array_4_io_d_in_0_b),
    .io_d_in_0_valid_b(array_4_io_d_in_0_valid_b),
    .io_d_in_1_a(array_4_io_d_in_1_a),
    .io_d_in_1_valid_a(array_4_io_d_in_1_valid_a),
    .io_d_in_1_b(array_4_io_d_in_1_b),
    .io_d_in_1_valid_b(array_4_io_d_in_1_valid_b),
    .io_d_in_2_a(array_4_io_d_in_2_a),
    .io_d_in_2_valid_a(array_4_io_d_in_2_valid_a),
    .io_d_in_2_b(array_4_io_d_in_2_b),
    .io_d_in_2_valid_b(array_4_io_d_in_2_valid_b),
    .io_d_in_3_a(array_4_io_d_in_3_a),
    .io_d_in_3_valid_a(array_4_io_d_in_3_valid_a),
    .io_d_in_3_b(array_4_io_d_in_3_b),
    .io_d_in_3_valid_b(array_4_io_d_in_3_valid_b),
    .io_d_in_4_a(array_4_io_d_in_4_a),
    .io_d_in_4_valid_a(array_4_io_d_in_4_valid_a),
    .io_d_in_4_b(array_4_io_d_in_4_b),
    .io_d_in_4_valid_b(array_4_io_d_in_4_valid_b),
    .io_d_in_5_a(array_4_io_d_in_5_a),
    .io_d_in_5_valid_a(array_4_io_d_in_5_valid_a),
    .io_d_in_5_b(array_4_io_d_in_5_b),
    .io_d_in_5_valid_b(array_4_io_d_in_5_valid_b),
    .io_d_in_6_a(array_4_io_d_in_6_a),
    .io_d_in_6_valid_a(array_4_io_d_in_6_valid_a),
    .io_d_in_6_b(array_4_io_d_in_6_b),
    .io_d_in_6_valid_b(array_4_io_d_in_6_valid_b),
    .io_d_in_7_a(array_4_io_d_in_7_a),
    .io_d_in_7_valid_a(array_4_io_d_in_7_valid_a),
    .io_d_in_7_b(array_4_io_d_in_7_b),
    .io_d_in_7_valid_b(array_4_io_d_in_7_valid_b),
    .io_d_in_8_a(array_4_io_d_in_8_a),
    .io_d_in_8_valid_a(array_4_io_d_in_8_valid_a),
    .io_d_in_8_b(array_4_io_d_in_8_b),
    .io_d_in_8_valid_b(array_4_io_d_in_8_valid_b),
    .io_d_in_9_a(array_4_io_d_in_9_a),
    .io_d_in_9_valid_a(array_4_io_d_in_9_valid_a),
    .io_d_in_9_b(array_4_io_d_in_9_b),
    .io_d_in_9_valid_b(array_4_io_d_in_9_valid_b),
    .io_d_in_10_a(array_4_io_d_in_10_a),
    .io_d_in_10_valid_a(array_4_io_d_in_10_valid_a),
    .io_d_in_10_b(array_4_io_d_in_10_b),
    .io_d_in_10_valid_b(array_4_io_d_in_10_valid_b),
    .io_d_in_11_a(array_4_io_d_in_11_a),
    .io_d_in_11_valid_a(array_4_io_d_in_11_valid_a),
    .io_d_in_11_b(array_4_io_d_in_11_b),
    .io_d_in_11_valid_b(array_4_io_d_in_11_valid_b),
    .io_d_in_12_a(array_4_io_d_in_12_a),
    .io_d_in_12_valid_a(array_4_io_d_in_12_valid_a),
    .io_d_in_12_b(array_4_io_d_in_12_b),
    .io_d_in_12_valid_b(array_4_io_d_in_12_valid_b),
    .io_d_in_13_a(array_4_io_d_in_13_a),
    .io_d_in_13_valid_a(array_4_io_d_in_13_valid_a),
    .io_d_in_13_b(array_4_io_d_in_13_b),
    .io_d_in_13_valid_b(array_4_io_d_in_13_valid_b),
    .io_d_in_14_a(array_4_io_d_in_14_a),
    .io_d_in_14_valid_a(array_4_io_d_in_14_valid_a),
    .io_d_in_14_b(array_4_io_d_in_14_b),
    .io_d_in_14_valid_b(array_4_io_d_in_14_valid_b),
    .io_d_in_15_a(array_4_io_d_in_15_a),
    .io_d_in_15_valid_a(array_4_io_d_in_15_valid_a),
    .io_d_in_15_b(array_4_io_d_in_15_b),
    .io_d_in_15_valid_b(array_4_io_d_in_15_valid_b),
    .io_d_in_16_a(array_4_io_d_in_16_a),
    .io_d_in_16_valid_a(array_4_io_d_in_16_valid_a),
    .io_d_in_16_b(array_4_io_d_in_16_b),
    .io_d_in_16_valid_b(array_4_io_d_in_16_valid_b),
    .io_d_in_17_a(array_4_io_d_in_17_a),
    .io_d_in_17_valid_a(array_4_io_d_in_17_valid_a),
    .io_d_in_17_b(array_4_io_d_in_17_b),
    .io_d_in_17_valid_b(array_4_io_d_in_17_valid_b),
    .io_d_in_18_a(array_4_io_d_in_18_a),
    .io_d_in_18_valid_a(array_4_io_d_in_18_valid_a),
    .io_d_in_18_b(array_4_io_d_in_18_b),
    .io_d_in_18_valid_b(array_4_io_d_in_18_valid_b),
    .io_d_in_19_a(array_4_io_d_in_19_a),
    .io_d_in_19_valid_a(array_4_io_d_in_19_valid_a),
    .io_d_in_19_b(array_4_io_d_in_19_b),
    .io_d_in_19_valid_b(array_4_io_d_in_19_valid_b),
    .io_d_in_20_a(array_4_io_d_in_20_a),
    .io_d_in_20_valid_a(array_4_io_d_in_20_valid_a),
    .io_d_in_20_b(array_4_io_d_in_20_b),
    .io_d_in_20_valid_b(array_4_io_d_in_20_valid_b),
    .io_d_in_21_a(array_4_io_d_in_21_a),
    .io_d_in_21_valid_a(array_4_io_d_in_21_valid_a),
    .io_d_in_21_b(array_4_io_d_in_21_b),
    .io_d_in_21_valid_b(array_4_io_d_in_21_valid_b),
    .io_d_in_22_a(array_4_io_d_in_22_a),
    .io_d_in_22_valid_a(array_4_io_d_in_22_valid_a),
    .io_d_in_22_b(array_4_io_d_in_22_b),
    .io_d_in_22_valid_b(array_4_io_d_in_22_valid_b),
    .io_d_in_23_a(array_4_io_d_in_23_a),
    .io_d_in_23_valid_a(array_4_io_d_in_23_valid_a),
    .io_d_in_23_b(array_4_io_d_in_23_b),
    .io_d_in_23_valid_b(array_4_io_d_in_23_valid_b),
    .io_d_in_24_a(array_4_io_d_in_24_a),
    .io_d_in_24_valid_a(array_4_io_d_in_24_valid_a),
    .io_d_in_24_b(array_4_io_d_in_24_b),
    .io_d_in_24_valid_b(array_4_io_d_in_24_valid_b),
    .io_d_in_25_a(array_4_io_d_in_25_a),
    .io_d_in_25_valid_a(array_4_io_d_in_25_valid_a),
    .io_d_in_25_b(array_4_io_d_in_25_b),
    .io_d_in_25_valid_b(array_4_io_d_in_25_valid_b),
    .io_d_in_26_a(array_4_io_d_in_26_a),
    .io_d_in_26_valid_a(array_4_io_d_in_26_valid_a),
    .io_d_in_26_b(array_4_io_d_in_26_b),
    .io_d_in_26_valid_b(array_4_io_d_in_26_valid_b),
    .io_d_in_27_a(array_4_io_d_in_27_a),
    .io_d_in_27_valid_a(array_4_io_d_in_27_valid_a),
    .io_d_in_27_b(array_4_io_d_in_27_b),
    .io_d_in_27_valid_b(array_4_io_d_in_27_valid_b),
    .io_d_in_28_a(array_4_io_d_in_28_a),
    .io_d_in_28_valid_a(array_4_io_d_in_28_valid_a),
    .io_d_in_28_b(array_4_io_d_in_28_b),
    .io_d_in_28_valid_b(array_4_io_d_in_28_valid_b),
    .io_d_in_29_a(array_4_io_d_in_29_a),
    .io_d_in_29_valid_a(array_4_io_d_in_29_valid_a),
    .io_d_in_29_b(array_4_io_d_in_29_b),
    .io_d_in_29_valid_b(array_4_io_d_in_29_valid_b),
    .io_d_in_30_a(array_4_io_d_in_30_a),
    .io_d_in_30_valid_a(array_4_io_d_in_30_valid_a),
    .io_d_in_30_b(array_4_io_d_in_30_b),
    .io_d_in_30_valid_b(array_4_io_d_in_30_valid_b),
    .io_d_in_31_a(array_4_io_d_in_31_a),
    .io_d_in_31_valid_a(array_4_io_d_in_31_valid_a),
    .io_d_in_31_b(array_4_io_d_in_31_b),
    .io_d_in_31_valid_b(array_4_io_d_in_31_valid_b),
    .io_d_out_0_a(array_4_io_d_out_0_a),
    .io_d_out_0_valid_a(array_4_io_d_out_0_valid_a),
    .io_d_out_0_b(array_4_io_d_out_0_b),
    .io_d_out_0_valid_b(array_4_io_d_out_0_valid_b),
    .io_d_out_1_a(array_4_io_d_out_1_a),
    .io_d_out_1_valid_a(array_4_io_d_out_1_valid_a),
    .io_d_out_1_b(array_4_io_d_out_1_b),
    .io_d_out_1_valid_b(array_4_io_d_out_1_valid_b),
    .io_d_out_2_a(array_4_io_d_out_2_a),
    .io_d_out_2_valid_a(array_4_io_d_out_2_valid_a),
    .io_d_out_2_b(array_4_io_d_out_2_b),
    .io_d_out_2_valid_b(array_4_io_d_out_2_valid_b),
    .io_d_out_3_a(array_4_io_d_out_3_a),
    .io_d_out_3_valid_a(array_4_io_d_out_3_valid_a),
    .io_d_out_3_b(array_4_io_d_out_3_b),
    .io_d_out_3_valid_b(array_4_io_d_out_3_valid_b),
    .io_d_out_4_a(array_4_io_d_out_4_a),
    .io_d_out_4_valid_a(array_4_io_d_out_4_valid_a),
    .io_d_out_4_b(array_4_io_d_out_4_b),
    .io_d_out_4_valid_b(array_4_io_d_out_4_valid_b),
    .io_d_out_5_a(array_4_io_d_out_5_a),
    .io_d_out_5_valid_a(array_4_io_d_out_5_valid_a),
    .io_d_out_5_b(array_4_io_d_out_5_b),
    .io_d_out_5_valid_b(array_4_io_d_out_5_valid_b),
    .io_d_out_6_a(array_4_io_d_out_6_a),
    .io_d_out_6_valid_a(array_4_io_d_out_6_valid_a),
    .io_d_out_6_b(array_4_io_d_out_6_b),
    .io_d_out_6_valid_b(array_4_io_d_out_6_valid_b),
    .io_d_out_7_a(array_4_io_d_out_7_a),
    .io_d_out_7_valid_a(array_4_io_d_out_7_valid_a),
    .io_d_out_7_b(array_4_io_d_out_7_b),
    .io_d_out_7_valid_b(array_4_io_d_out_7_valid_b),
    .io_d_out_8_a(array_4_io_d_out_8_a),
    .io_d_out_8_valid_a(array_4_io_d_out_8_valid_a),
    .io_d_out_8_b(array_4_io_d_out_8_b),
    .io_d_out_8_valid_b(array_4_io_d_out_8_valid_b),
    .io_d_out_9_a(array_4_io_d_out_9_a),
    .io_d_out_9_valid_a(array_4_io_d_out_9_valid_a),
    .io_d_out_9_b(array_4_io_d_out_9_b),
    .io_d_out_9_valid_b(array_4_io_d_out_9_valid_b),
    .io_d_out_10_a(array_4_io_d_out_10_a),
    .io_d_out_10_valid_a(array_4_io_d_out_10_valid_a),
    .io_d_out_10_b(array_4_io_d_out_10_b),
    .io_d_out_10_valid_b(array_4_io_d_out_10_valid_b),
    .io_d_out_11_a(array_4_io_d_out_11_a),
    .io_d_out_11_valid_a(array_4_io_d_out_11_valid_a),
    .io_d_out_11_b(array_4_io_d_out_11_b),
    .io_d_out_11_valid_b(array_4_io_d_out_11_valid_b),
    .io_d_out_12_a(array_4_io_d_out_12_a),
    .io_d_out_12_valid_a(array_4_io_d_out_12_valid_a),
    .io_d_out_12_b(array_4_io_d_out_12_b),
    .io_d_out_12_valid_b(array_4_io_d_out_12_valid_b),
    .io_d_out_13_a(array_4_io_d_out_13_a),
    .io_d_out_13_valid_a(array_4_io_d_out_13_valid_a),
    .io_d_out_13_b(array_4_io_d_out_13_b),
    .io_d_out_13_valid_b(array_4_io_d_out_13_valid_b),
    .io_d_out_14_a(array_4_io_d_out_14_a),
    .io_d_out_14_valid_a(array_4_io_d_out_14_valid_a),
    .io_d_out_14_b(array_4_io_d_out_14_b),
    .io_d_out_14_valid_b(array_4_io_d_out_14_valid_b),
    .io_d_out_15_a(array_4_io_d_out_15_a),
    .io_d_out_15_valid_a(array_4_io_d_out_15_valid_a),
    .io_d_out_15_b(array_4_io_d_out_15_b),
    .io_d_out_15_valid_b(array_4_io_d_out_15_valid_b),
    .io_d_out_16_a(array_4_io_d_out_16_a),
    .io_d_out_16_valid_a(array_4_io_d_out_16_valid_a),
    .io_d_out_16_b(array_4_io_d_out_16_b),
    .io_d_out_16_valid_b(array_4_io_d_out_16_valid_b),
    .io_d_out_17_a(array_4_io_d_out_17_a),
    .io_d_out_17_valid_a(array_4_io_d_out_17_valid_a),
    .io_d_out_17_b(array_4_io_d_out_17_b),
    .io_d_out_17_valid_b(array_4_io_d_out_17_valid_b),
    .io_d_out_18_a(array_4_io_d_out_18_a),
    .io_d_out_18_valid_a(array_4_io_d_out_18_valid_a),
    .io_d_out_18_b(array_4_io_d_out_18_b),
    .io_d_out_18_valid_b(array_4_io_d_out_18_valid_b),
    .io_d_out_19_a(array_4_io_d_out_19_a),
    .io_d_out_19_valid_a(array_4_io_d_out_19_valid_a),
    .io_d_out_19_b(array_4_io_d_out_19_b),
    .io_d_out_19_valid_b(array_4_io_d_out_19_valid_b),
    .io_d_out_20_a(array_4_io_d_out_20_a),
    .io_d_out_20_valid_a(array_4_io_d_out_20_valid_a),
    .io_d_out_20_b(array_4_io_d_out_20_b),
    .io_d_out_20_valid_b(array_4_io_d_out_20_valid_b),
    .io_d_out_21_a(array_4_io_d_out_21_a),
    .io_d_out_21_valid_a(array_4_io_d_out_21_valid_a),
    .io_d_out_21_b(array_4_io_d_out_21_b),
    .io_d_out_21_valid_b(array_4_io_d_out_21_valid_b),
    .io_d_out_22_a(array_4_io_d_out_22_a),
    .io_d_out_22_valid_a(array_4_io_d_out_22_valid_a),
    .io_d_out_22_b(array_4_io_d_out_22_b),
    .io_d_out_22_valid_b(array_4_io_d_out_22_valid_b),
    .io_d_out_23_a(array_4_io_d_out_23_a),
    .io_d_out_23_valid_a(array_4_io_d_out_23_valid_a),
    .io_d_out_23_b(array_4_io_d_out_23_b),
    .io_d_out_23_valid_b(array_4_io_d_out_23_valid_b),
    .io_d_out_24_a(array_4_io_d_out_24_a),
    .io_d_out_24_valid_a(array_4_io_d_out_24_valid_a),
    .io_d_out_24_b(array_4_io_d_out_24_b),
    .io_d_out_24_valid_b(array_4_io_d_out_24_valid_b),
    .io_d_out_25_a(array_4_io_d_out_25_a),
    .io_d_out_25_valid_a(array_4_io_d_out_25_valid_a),
    .io_d_out_25_b(array_4_io_d_out_25_b),
    .io_d_out_25_valid_b(array_4_io_d_out_25_valid_b),
    .io_d_out_26_a(array_4_io_d_out_26_a),
    .io_d_out_26_valid_a(array_4_io_d_out_26_valid_a),
    .io_d_out_26_b(array_4_io_d_out_26_b),
    .io_d_out_26_valid_b(array_4_io_d_out_26_valid_b),
    .io_d_out_27_a(array_4_io_d_out_27_a),
    .io_d_out_27_valid_a(array_4_io_d_out_27_valid_a),
    .io_d_out_27_b(array_4_io_d_out_27_b),
    .io_d_out_27_valid_b(array_4_io_d_out_27_valid_b),
    .io_d_out_28_a(array_4_io_d_out_28_a),
    .io_d_out_28_valid_a(array_4_io_d_out_28_valid_a),
    .io_d_out_28_b(array_4_io_d_out_28_b),
    .io_d_out_28_valid_b(array_4_io_d_out_28_valid_b),
    .io_d_out_29_a(array_4_io_d_out_29_a),
    .io_d_out_29_valid_a(array_4_io_d_out_29_valid_a),
    .io_d_out_29_b(array_4_io_d_out_29_b),
    .io_d_out_29_valid_b(array_4_io_d_out_29_valid_b),
    .io_d_out_30_a(array_4_io_d_out_30_a),
    .io_d_out_30_valid_a(array_4_io_d_out_30_valid_a),
    .io_d_out_30_b(array_4_io_d_out_30_b),
    .io_d_out_30_valid_b(array_4_io_d_out_30_valid_b),
    .io_d_out_31_a(array_4_io_d_out_31_a),
    .io_d_out_31_valid_a(array_4_io_d_out_31_valid_a),
    .io_d_out_31_b(array_4_io_d_out_31_b),
    .io_d_out_31_valid_b(array_4_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_4_io_wr_en_mem1),
    .io_wr_en_mem2(array_4_io_wr_en_mem2),
    .io_wr_en_mem3(array_4_io_wr_en_mem3),
    .io_wr_en_mem4(array_4_io_wr_en_mem4),
    .io_wr_en_mem5(array_4_io_wr_en_mem5),
    .io_wr_en_mem6(array_4_io_wr_en_mem6),
    .io_wr_instr_mem1(array_4_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_4_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_4_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_4_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_4_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_4_io_wr_instr_mem6),
    .io_PC1_in(array_4_io_PC1_in),
    .io_PC6_out(array_4_io_PC6_out),
    .io_Addr_in(array_4_io_Addr_in),
    .io_Addr_out(array_4_io_Addr_out)
  );
  BuildingBlockNew array_5 ( // @[BP.scala 45:51]
    .clock(array_5_clock),
    .reset(array_5_reset),
    .io_d_in_0_a(array_5_io_d_in_0_a),
    .io_d_in_0_valid_a(array_5_io_d_in_0_valid_a),
    .io_d_in_0_b(array_5_io_d_in_0_b),
    .io_d_in_0_valid_b(array_5_io_d_in_0_valid_b),
    .io_d_in_1_a(array_5_io_d_in_1_a),
    .io_d_in_1_valid_a(array_5_io_d_in_1_valid_a),
    .io_d_in_1_b(array_5_io_d_in_1_b),
    .io_d_in_1_valid_b(array_5_io_d_in_1_valid_b),
    .io_d_in_2_a(array_5_io_d_in_2_a),
    .io_d_in_2_valid_a(array_5_io_d_in_2_valid_a),
    .io_d_in_2_b(array_5_io_d_in_2_b),
    .io_d_in_2_valid_b(array_5_io_d_in_2_valid_b),
    .io_d_in_3_a(array_5_io_d_in_3_a),
    .io_d_in_3_valid_a(array_5_io_d_in_3_valid_a),
    .io_d_in_3_b(array_5_io_d_in_3_b),
    .io_d_in_3_valid_b(array_5_io_d_in_3_valid_b),
    .io_d_in_4_a(array_5_io_d_in_4_a),
    .io_d_in_4_valid_a(array_5_io_d_in_4_valid_a),
    .io_d_in_4_b(array_5_io_d_in_4_b),
    .io_d_in_4_valid_b(array_5_io_d_in_4_valid_b),
    .io_d_in_5_a(array_5_io_d_in_5_a),
    .io_d_in_5_valid_a(array_5_io_d_in_5_valid_a),
    .io_d_in_5_b(array_5_io_d_in_5_b),
    .io_d_in_5_valid_b(array_5_io_d_in_5_valid_b),
    .io_d_in_6_a(array_5_io_d_in_6_a),
    .io_d_in_6_valid_a(array_5_io_d_in_6_valid_a),
    .io_d_in_6_b(array_5_io_d_in_6_b),
    .io_d_in_6_valid_b(array_5_io_d_in_6_valid_b),
    .io_d_in_7_a(array_5_io_d_in_7_a),
    .io_d_in_7_valid_a(array_5_io_d_in_7_valid_a),
    .io_d_in_7_b(array_5_io_d_in_7_b),
    .io_d_in_7_valid_b(array_5_io_d_in_7_valid_b),
    .io_d_in_8_a(array_5_io_d_in_8_a),
    .io_d_in_8_valid_a(array_5_io_d_in_8_valid_a),
    .io_d_in_8_b(array_5_io_d_in_8_b),
    .io_d_in_8_valid_b(array_5_io_d_in_8_valid_b),
    .io_d_in_9_a(array_5_io_d_in_9_a),
    .io_d_in_9_valid_a(array_5_io_d_in_9_valid_a),
    .io_d_in_9_b(array_5_io_d_in_9_b),
    .io_d_in_9_valid_b(array_5_io_d_in_9_valid_b),
    .io_d_in_10_a(array_5_io_d_in_10_a),
    .io_d_in_10_valid_a(array_5_io_d_in_10_valid_a),
    .io_d_in_10_b(array_5_io_d_in_10_b),
    .io_d_in_10_valid_b(array_5_io_d_in_10_valid_b),
    .io_d_in_11_a(array_5_io_d_in_11_a),
    .io_d_in_11_valid_a(array_5_io_d_in_11_valid_a),
    .io_d_in_11_b(array_5_io_d_in_11_b),
    .io_d_in_11_valid_b(array_5_io_d_in_11_valid_b),
    .io_d_in_12_a(array_5_io_d_in_12_a),
    .io_d_in_12_valid_a(array_5_io_d_in_12_valid_a),
    .io_d_in_12_b(array_5_io_d_in_12_b),
    .io_d_in_12_valid_b(array_5_io_d_in_12_valid_b),
    .io_d_in_13_a(array_5_io_d_in_13_a),
    .io_d_in_13_valid_a(array_5_io_d_in_13_valid_a),
    .io_d_in_13_b(array_5_io_d_in_13_b),
    .io_d_in_13_valid_b(array_5_io_d_in_13_valid_b),
    .io_d_in_14_a(array_5_io_d_in_14_a),
    .io_d_in_14_valid_a(array_5_io_d_in_14_valid_a),
    .io_d_in_14_b(array_5_io_d_in_14_b),
    .io_d_in_14_valid_b(array_5_io_d_in_14_valid_b),
    .io_d_in_15_a(array_5_io_d_in_15_a),
    .io_d_in_15_valid_a(array_5_io_d_in_15_valid_a),
    .io_d_in_15_b(array_5_io_d_in_15_b),
    .io_d_in_15_valid_b(array_5_io_d_in_15_valid_b),
    .io_d_in_16_a(array_5_io_d_in_16_a),
    .io_d_in_16_valid_a(array_5_io_d_in_16_valid_a),
    .io_d_in_16_b(array_5_io_d_in_16_b),
    .io_d_in_16_valid_b(array_5_io_d_in_16_valid_b),
    .io_d_in_17_a(array_5_io_d_in_17_a),
    .io_d_in_17_valid_a(array_5_io_d_in_17_valid_a),
    .io_d_in_17_b(array_5_io_d_in_17_b),
    .io_d_in_17_valid_b(array_5_io_d_in_17_valid_b),
    .io_d_in_18_a(array_5_io_d_in_18_a),
    .io_d_in_18_valid_a(array_5_io_d_in_18_valid_a),
    .io_d_in_18_b(array_5_io_d_in_18_b),
    .io_d_in_18_valid_b(array_5_io_d_in_18_valid_b),
    .io_d_in_19_a(array_5_io_d_in_19_a),
    .io_d_in_19_valid_a(array_5_io_d_in_19_valid_a),
    .io_d_in_19_b(array_5_io_d_in_19_b),
    .io_d_in_19_valid_b(array_5_io_d_in_19_valid_b),
    .io_d_in_20_a(array_5_io_d_in_20_a),
    .io_d_in_20_valid_a(array_5_io_d_in_20_valid_a),
    .io_d_in_20_b(array_5_io_d_in_20_b),
    .io_d_in_20_valid_b(array_5_io_d_in_20_valid_b),
    .io_d_in_21_a(array_5_io_d_in_21_a),
    .io_d_in_21_valid_a(array_5_io_d_in_21_valid_a),
    .io_d_in_21_b(array_5_io_d_in_21_b),
    .io_d_in_21_valid_b(array_5_io_d_in_21_valid_b),
    .io_d_in_22_a(array_5_io_d_in_22_a),
    .io_d_in_22_valid_a(array_5_io_d_in_22_valid_a),
    .io_d_in_22_b(array_5_io_d_in_22_b),
    .io_d_in_22_valid_b(array_5_io_d_in_22_valid_b),
    .io_d_in_23_a(array_5_io_d_in_23_a),
    .io_d_in_23_valid_a(array_5_io_d_in_23_valid_a),
    .io_d_in_23_b(array_5_io_d_in_23_b),
    .io_d_in_23_valid_b(array_5_io_d_in_23_valid_b),
    .io_d_in_24_a(array_5_io_d_in_24_a),
    .io_d_in_24_valid_a(array_5_io_d_in_24_valid_a),
    .io_d_in_24_b(array_5_io_d_in_24_b),
    .io_d_in_24_valid_b(array_5_io_d_in_24_valid_b),
    .io_d_in_25_a(array_5_io_d_in_25_a),
    .io_d_in_25_valid_a(array_5_io_d_in_25_valid_a),
    .io_d_in_25_b(array_5_io_d_in_25_b),
    .io_d_in_25_valid_b(array_5_io_d_in_25_valid_b),
    .io_d_in_26_a(array_5_io_d_in_26_a),
    .io_d_in_26_valid_a(array_5_io_d_in_26_valid_a),
    .io_d_in_26_b(array_5_io_d_in_26_b),
    .io_d_in_26_valid_b(array_5_io_d_in_26_valid_b),
    .io_d_in_27_a(array_5_io_d_in_27_a),
    .io_d_in_27_valid_a(array_5_io_d_in_27_valid_a),
    .io_d_in_27_b(array_5_io_d_in_27_b),
    .io_d_in_27_valid_b(array_5_io_d_in_27_valid_b),
    .io_d_in_28_a(array_5_io_d_in_28_a),
    .io_d_in_28_valid_a(array_5_io_d_in_28_valid_a),
    .io_d_in_28_b(array_5_io_d_in_28_b),
    .io_d_in_28_valid_b(array_5_io_d_in_28_valid_b),
    .io_d_in_29_a(array_5_io_d_in_29_a),
    .io_d_in_29_valid_a(array_5_io_d_in_29_valid_a),
    .io_d_in_29_b(array_5_io_d_in_29_b),
    .io_d_in_29_valid_b(array_5_io_d_in_29_valid_b),
    .io_d_in_30_a(array_5_io_d_in_30_a),
    .io_d_in_30_valid_a(array_5_io_d_in_30_valid_a),
    .io_d_in_30_b(array_5_io_d_in_30_b),
    .io_d_in_30_valid_b(array_5_io_d_in_30_valid_b),
    .io_d_in_31_a(array_5_io_d_in_31_a),
    .io_d_in_31_valid_a(array_5_io_d_in_31_valid_a),
    .io_d_in_31_b(array_5_io_d_in_31_b),
    .io_d_in_31_valid_b(array_5_io_d_in_31_valid_b),
    .io_d_out_0_a(array_5_io_d_out_0_a),
    .io_d_out_0_valid_a(array_5_io_d_out_0_valid_a),
    .io_d_out_0_b(array_5_io_d_out_0_b),
    .io_d_out_0_valid_b(array_5_io_d_out_0_valid_b),
    .io_d_out_1_a(array_5_io_d_out_1_a),
    .io_d_out_1_valid_a(array_5_io_d_out_1_valid_a),
    .io_d_out_1_b(array_5_io_d_out_1_b),
    .io_d_out_1_valid_b(array_5_io_d_out_1_valid_b),
    .io_d_out_2_a(array_5_io_d_out_2_a),
    .io_d_out_2_valid_a(array_5_io_d_out_2_valid_a),
    .io_d_out_2_b(array_5_io_d_out_2_b),
    .io_d_out_2_valid_b(array_5_io_d_out_2_valid_b),
    .io_d_out_3_a(array_5_io_d_out_3_a),
    .io_d_out_3_valid_a(array_5_io_d_out_3_valid_a),
    .io_d_out_3_b(array_5_io_d_out_3_b),
    .io_d_out_3_valid_b(array_5_io_d_out_3_valid_b),
    .io_d_out_4_a(array_5_io_d_out_4_a),
    .io_d_out_4_valid_a(array_5_io_d_out_4_valid_a),
    .io_d_out_4_b(array_5_io_d_out_4_b),
    .io_d_out_4_valid_b(array_5_io_d_out_4_valid_b),
    .io_d_out_5_a(array_5_io_d_out_5_a),
    .io_d_out_5_valid_a(array_5_io_d_out_5_valid_a),
    .io_d_out_5_b(array_5_io_d_out_5_b),
    .io_d_out_5_valid_b(array_5_io_d_out_5_valid_b),
    .io_d_out_6_a(array_5_io_d_out_6_a),
    .io_d_out_6_valid_a(array_5_io_d_out_6_valid_a),
    .io_d_out_6_b(array_5_io_d_out_6_b),
    .io_d_out_6_valid_b(array_5_io_d_out_6_valid_b),
    .io_d_out_7_a(array_5_io_d_out_7_a),
    .io_d_out_7_valid_a(array_5_io_d_out_7_valid_a),
    .io_d_out_7_b(array_5_io_d_out_7_b),
    .io_d_out_7_valid_b(array_5_io_d_out_7_valid_b),
    .io_d_out_8_a(array_5_io_d_out_8_a),
    .io_d_out_8_valid_a(array_5_io_d_out_8_valid_a),
    .io_d_out_8_b(array_5_io_d_out_8_b),
    .io_d_out_8_valid_b(array_5_io_d_out_8_valid_b),
    .io_d_out_9_a(array_5_io_d_out_9_a),
    .io_d_out_9_valid_a(array_5_io_d_out_9_valid_a),
    .io_d_out_9_b(array_5_io_d_out_9_b),
    .io_d_out_9_valid_b(array_5_io_d_out_9_valid_b),
    .io_d_out_10_a(array_5_io_d_out_10_a),
    .io_d_out_10_valid_a(array_5_io_d_out_10_valid_a),
    .io_d_out_10_b(array_5_io_d_out_10_b),
    .io_d_out_10_valid_b(array_5_io_d_out_10_valid_b),
    .io_d_out_11_a(array_5_io_d_out_11_a),
    .io_d_out_11_valid_a(array_5_io_d_out_11_valid_a),
    .io_d_out_11_b(array_5_io_d_out_11_b),
    .io_d_out_11_valid_b(array_5_io_d_out_11_valid_b),
    .io_d_out_12_a(array_5_io_d_out_12_a),
    .io_d_out_12_valid_a(array_5_io_d_out_12_valid_a),
    .io_d_out_12_b(array_5_io_d_out_12_b),
    .io_d_out_12_valid_b(array_5_io_d_out_12_valid_b),
    .io_d_out_13_a(array_5_io_d_out_13_a),
    .io_d_out_13_valid_a(array_5_io_d_out_13_valid_a),
    .io_d_out_13_b(array_5_io_d_out_13_b),
    .io_d_out_13_valid_b(array_5_io_d_out_13_valid_b),
    .io_d_out_14_a(array_5_io_d_out_14_a),
    .io_d_out_14_valid_a(array_5_io_d_out_14_valid_a),
    .io_d_out_14_b(array_5_io_d_out_14_b),
    .io_d_out_14_valid_b(array_5_io_d_out_14_valid_b),
    .io_d_out_15_a(array_5_io_d_out_15_a),
    .io_d_out_15_valid_a(array_5_io_d_out_15_valid_a),
    .io_d_out_15_b(array_5_io_d_out_15_b),
    .io_d_out_15_valid_b(array_5_io_d_out_15_valid_b),
    .io_d_out_16_a(array_5_io_d_out_16_a),
    .io_d_out_16_valid_a(array_5_io_d_out_16_valid_a),
    .io_d_out_16_b(array_5_io_d_out_16_b),
    .io_d_out_16_valid_b(array_5_io_d_out_16_valid_b),
    .io_d_out_17_a(array_5_io_d_out_17_a),
    .io_d_out_17_valid_a(array_5_io_d_out_17_valid_a),
    .io_d_out_17_b(array_5_io_d_out_17_b),
    .io_d_out_17_valid_b(array_5_io_d_out_17_valid_b),
    .io_d_out_18_a(array_5_io_d_out_18_a),
    .io_d_out_18_valid_a(array_5_io_d_out_18_valid_a),
    .io_d_out_18_b(array_5_io_d_out_18_b),
    .io_d_out_18_valid_b(array_5_io_d_out_18_valid_b),
    .io_d_out_19_a(array_5_io_d_out_19_a),
    .io_d_out_19_valid_a(array_5_io_d_out_19_valid_a),
    .io_d_out_19_b(array_5_io_d_out_19_b),
    .io_d_out_19_valid_b(array_5_io_d_out_19_valid_b),
    .io_d_out_20_a(array_5_io_d_out_20_a),
    .io_d_out_20_valid_a(array_5_io_d_out_20_valid_a),
    .io_d_out_20_b(array_5_io_d_out_20_b),
    .io_d_out_20_valid_b(array_5_io_d_out_20_valid_b),
    .io_d_out_21_a(array_5_io_d_out_21_a),
    .io_d_out_21_valid_a(array_5_io_d_out_21_valid_a),
    .io_d_out_21_b(array_5_io_d_out_21_b),
    .io_d_out_21_valid_b(array_5_io_d_out_21_valid_b),
    .io_d_out_22_a(array_5_io_d_out_22_a),
    .io_d_out_22_valid_a(array_5_io_d_out_22_valid_a),
    .io_d_out_22_b(array_5_io_d_out_22_b),
    .io_d_out_22_valid_b(array_5_io_d_out_22_valid_b),
    .io_d_out_23_a(array_5_io_d_out_23_a),
    .io_d_out_23_valid_a(array_5_io_d_out_23_valid_a),
    .io_d_out_23_b(array_5_io_d_out_23_b),
    .io_d_out_23_valid_b(array_5_io_d_out_23_valid_b),
    .io_d_out_24_a(array_5_io_d_out_24_a),
    .io_d_out_24_valid_a(array_5_io_d_out_24_valid_a),
    .io_d_out_24_b(array_5_io_d_out_24_b),
    .io_d_out_24_valid_b(array_5_io_d_out_24_valid_b),
    .io_d_out_25_a(array_5_io_d_out_25_a),
    .io_d_out_25_valid_a(array_5_io_d_out_25_valid_a),
    .io_d_out_25_b(array_5_io_d_out_25_b),
    .io_d_out_25_valid_b(array_5_io_d_out_25_valid_b),
    .io_d_out_26_a(array_5_io_d_out_26_a),
    .io_d_out_26_valid_a(array_5_io_d_out_26_valid_a),
    .io_d_out_26_b(array_5_io_d_out_26_b),
    .io_d_out_26_valid_b(array_5_io_d_out_26_valid_b),
    .io_d_out_27_a(array_5_io_d_out_27_a),
    .io_d_out_27_valid_a(array_5_io_d_out_27_valid_a),
    .io_d_out_27_b(array_5_io_d_out_27_b),
    .io_d_out_27_valid_b(array_5_io_d_out_27_valid_b),
    .io_d_out_28_a(array_5_io_d_out_28_a),
    .io_d_out_28_valid_a(array_5_io_d_out_28_valid_a),
    .io_d_out_28_b(array_5_io_d_out_28_b),
    .io_d_out_28_valid_b(array_5_io_d_out_28_valid_b),
    .io_d_out_29_a(array_5_io_d_out_29_a),
    .io_d_out_29_valid_a(array_5_io_d_out_29_valid_a),
    .io_d_out_29_b(array_5_io_d_out_29_b),
    .io_d_out_29_valid_b(array_5_io_d_out_29_valid_b),
    .io_d_out_30_a(array_5_io_d_out_30_a),
    .io_d_out_30_valid_a(array_5_io_d_out_30_valid_a),
    .io_d_out_30_b(array_5_io_d_out_30_b),
    .io_d_out_30_valid_b(array_5_io_d_out_30_valid_b),
    .io_d_out_31_a(array_5_io_d_out_31_a),
    .io_d_out_31_valid_a(array_5_io_d_out_31_valid_a),
    .io_d_out_31_b(array_5_io_d_out_31_b),
    .io_d_out_31_valid_b(array_5_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_5_io_wr_en_mem1),
    .io_wr_en_mem2(array_5_io_wr_en_mem2),
    .io_wr_en_mem3(array_5_io_wr_en_mem3),
    .io_wr_en_mem4(array_5_io_wr_en_mem4),
    .io_wr_en_mem5(array_5_io_wr_en_mem5),
    .io_wr_en_mem6(array_5_io_wr_en_mem6),
    .io_wr_instr_mem1(array_5_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_5_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_5_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_5_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_5_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_5_io_wr_instr_mem6),
    .io_PC1_in(array_5_io_PC1_in),
    .io_PC6_out(array_5_io_PC6_out),
    .io_Addr_in(array_5_io_Addr_in),
    .io_Addr_out(array_5_io_Addr_out)
  );
  BuildingBlockNew array_6 ( // @[BP.scala 45:51]
    .clock(array_6_clock),
    .reset(array_6_reset),
    .io_d_in_0_a(array_6_io_d_in_0_a),
    .io_d_in_0_valid_a(array_6_io_d_in_0_valid_a),
    .io_d_in_0_b(array_6_io_d_in_0_b),
    .io_d_in_0_valid_b(array_6_io_d_in_0_valid_b),
    .io_d_in_1_a(array_6_io_d_in_1_a),
    .io_d_in_1_valid_a(array_6_io_d_in_1_valid_a),
    .io_d_in_1_b(array_6_io_d_in_1_b),
    .io_d_in_1_valid_b(array_6_io_d_in_1_valid_b),
    .io_d_in_2_a(array_6_io_d_in_2_a),
    .io_d_in_2_valid_a(array_6_io_d_in_2_valid_a),
    .io_d_in_2_b(array_6_io_d_in_2_b),
    .io_d_in_2_valid_b(array_6_io_d_in_2_valid_b),
    .io_d_in_3_a(array_6_io_d_in_3_a),
    .io_d_in_3_valid_a(array_6_io_d_in_3_valid_a),
    .io_d_in_3_b(array_6_io_d_in_3_b),
    .io_d_in_3_valid_b(array_6_io_d_in_3_valid_b),
    .io_d_in_4_a(array_6_io_d_in_4_a),
    .io_d_in_4_valid_a(array_6_io_d_in_4_valid_a),
    .io_d_in_4_b(array_6_io_d_in_4_b),
    .io_d_in_4_valid_b(array_6_io_d_in_4_valid_b),
    .io_d_in_5_a(array_6_io_d_in_5_a),
    .io_d_in_5_valid_a(array_6_io_d_in_5_valid_a),
    .io_d_in_5_b(array_6_io_d_in_5_b),
    .io_d_in_5_valid_b(array_6_io_d_in_5_valid_b),
    .io_d_in_6_a(array_6_io_d_in_6_a),
    .io_d_in_6_valid_a(array_6_io_d_in_6_valid_a),
    .io_d_in_6_b(array_6_io_d_in_6_b),
    .io_d_in_6_valid_b(array_6_io_d_in_6_valid_b),
    .io_d_in_7_a(array_6_io_d_in_7_a),
    .io_d_in_7_valid_a(array_6_io_d_in_7_valid_a),
    .io_d_in_7_b(array_6_io_d_in_7_b),
    .io_d_in_7_valid_b(array_6_io_d_in_7_valid_b),
    .io_d_in_8_a(array_6_io_d_in_8_a),
    .io_d_in_8_valid_a(array_6_io_d_in_8_valid_a),
    .io_d_in_8_b(array_6_io_d_in_8_b),
    .io_d_in_8_valid_b(array_6_io_d_in_8_valid_b),
    .io_d_in_9_a(array_6_io_d_in_9_a),
    .io_d_in_9_valid_a(array_6_io_d_in_9_valid_a),
    .io_d_in_9_b(array_6_io_d_in_9_b),
    .io_d_in_9_valid_b(array_6_io_d_in_9_valid_b),
    .io_d_in_10_a(array_6_io_d_in_10_a),
    .io_d_in_10_valid_a(array_6_io_d_in_10_valid_a),
    .io_d_in_10_b(array_6_io_d_in_10_b),
    .io_d_in_10_valid_b(array_6_io_d_in_10_valid_b),
    .io_d_in_11_a(array_6_io_d_in_11_a),
    .io_d_in_11_valid_a(array_6_io_d_in_11_valid_a),
    .io_d_in_11_b(array_6_io_d_in_11_b),
    .io_d_in_11_valid_b(array_6_io_d_in_11_valid_b),
    .io_d_in_12_a(array_6_io_d_in_12_a),
    .io_d_in_12_valid_a(array_6_io_d_in_12_valid_a),
    .io_d_in_12_b(array_6_io_d_in_12_b),
    .io_d_in_12_valid_b(array_6_io_d_in_12_valid_b),
    .io_d_in_13_a(array_6_io_d_in_13_a),
    .io_d_in_13_valid_a(array_6_io_d_in_13_valid_a),
    .io_d_in_13_b(array_6_io_d_in_13_b),
    .io_d_in_13_valid_b(array_6_io_d_in_13_valid_b),
    .io_d_in_14_a(array_6_io_d_in_14_a),
    .io_d_in_14_valid_a(array_6_io_d_in_14_valid_a),
    .io_d_in_14_b(array_6_io_d_in_14_b),
    .io_d_in_14_valid_b(array_6_io_d_in_14_valid_b),
    .io_d_in_15_a(array_6_io_d_in_15_a),
    .io_d_in_15_valid_a(array_6_io_d_in_15_valid_a),
    .io_d_in_15_b(array_6_io_d_in_15_b),
    .io_d_in_15_valid_b(array_6_io_d_in_15_valid_b),
    .io_d_in_16_a(array_6_io_d_in_16_a),
    .io_d_in_16_valid_a(array_6_io_d_in_16_valid_a),
    .io_d_in_16_b(array_6_io_d_in_16_b),
    .io_d_in_16_valid_b(array_6_io_d_in_16_valid_b),
    .io_d_in_17_a(array_6_io_d_in_17_a),
    .io_d_in_17_valid_a(array_6_io_d_in_17_valid_a),
    .io_d_in_17_b(array_6_io_d_in_17_b),
    .io_d_in_17_valid_b(array_6_io_d_in_17_valid_b),
    .io_d_in_18_a(array_6_io_d_in_18_a),
    .io_d_in_18_valid_a(array_6_io_d_in_18_valid_a),
    .io_d_in_18_b(array_6_io_d_in_18_b),
    .io_d_in_18_valid_b(array_6_io_d_in_18_valid_b),
    .io_d_in_19_a(array_6_io_d_in_19_a),
    .io_d_in_19_valid_a(array_6_io_d_in_19_valid_a),
    .io_d_in_19_b(array_6_io_d_in_19_b),
    .io_d_in_19_valid_b(array_6_io_d_in_19_valid_b),
    .io_d_in_20_a(array_6_io_d_in_20_a),
    .io_d_in_20_valid_a(array_6_io_d_in_20_valid_a),
    .io_d_in_20_b(array_6_io_d_in_20_b),
    .io_d_in_20_valid_b(array_6_io_d_in_20_valid_b),
    .io_d_in_21_a(array_6_io_d_in_21_a),
    .io_d_in_21_valid_a(array_6_io_d_in_21_valid_a),
    .io_d_in_21_b(array_6_io_d_in_21_b),
    .io_d_in_21_valid_b(array_6_io_d_in_21_valid_b),
    .io_d_in_22_a(array_6_io_d_in_22_a),
    .io_d_in_22_valid_a(array_6_io_d_in_22_valid_a),
    .io_d_in_22_b(array_6_io_d_in_22_b),
    .io_d_in_22_valid_b(array_6_io_d_in_22_valid_b),
    .io_d_in_23_a(array_6_io_d_in_23_a),
    .io_d_in_23_valid_a(array_6_io_d_in_23_valid_a),
    .io_d_in_23_b(array_6_io_d_in_23_b),
    .io_d_in_23_valid_b(array_6_io_d_in_23_valid_b),
    .io_d_in_24_a(array_6_io_d_in_24_a),
    .io_d_in_24_valid_a(array_6_io_d_in_24_valid_a),
    .io_d_in_24_b(array_6_io_d_in_24_b),
    .io_d_in_24_valid_b(array_6_io_d_in_24_valid_b),
    .io_d_in_25_a(array_6_io_d_in_25_a),
    .io_d_in_25_valid_a(array_6_io_d_in_25_valid_a),
    .io_d_in_25_b(array_6_io_d_in_25_b),
    .io_d_in_25_valid_b(array_6_io_d_in_25_valid_b),
    .io_d_in_26_a(array_6_io_d_in_26_a),
    .io_d_in_26_valid_a(array_6_io_d_in_26_valid_a),
    .io_d_in_26_b(array_6_io_d_in_26_b),
    .io_d_in_26_valid_b(array_6_io_d_in_26_valid_b),
    .io_d_in_27_a(array_6_io_d_in_27_a),
    .io_d_in_27_valid_a(array_6_io_d_in_27_valid_a),
    .io_d_in_27_b(array_6_io_d_in_27_b),
    .io_d_in_27_valid_b(array_6_io_d_in_27_valid_b),
    .io_d_in_28_a(array_6_io_d_in_28_a),
    .io_d_in_28_valid_a(array_6_io_d_in_28_valid_a),
    .io_d_in_28_b(array_6_io_d_in_28_b),
    .io_d_in_28_valid_b(array_6_io_d_in_28_valid_b),
    .io_d_in_29_a(array_6_io_d_in_29_a),
    .io_d_in_29_valid_a(array_6_io_d_in_29_valid_a),
    .io_d_in_29_b(array_6_io_d_in_29_b),
    .io_d_in_29_valid_b(array_6_io_d_in_29_valid_b),
    .io_d_in_30_a(array_6_io_d_in_30_a),
    .io_d_in_30_valid_a(array_6_io_d_in_30_valid_a),
    .io_d_in_30_b(array_6_io_d_in_30_b),
    .io_d_in_30_valid_b(array_6_io_d_in_30_valid_b),
    .io_d_in_31_a(array_6_io_d_in_31_a),
    .io_d_in_31_valid_a(array_6_io_d_in_31_valid_a),
    .io_d_in_31_b(array_6_io_d_in_31_b),
    .io_d_in_31_valid_b(array_6_io_d_in_31_valid_b),
    .io_d_out_0_a(array_6_io_d_out_0_a),
    .io_d_out_0_valid_a(array_6_io_d_out_0_valid_a),
    .io_d_out_0_b(array_6_io_d_out_0_b),
    .io_d_out_0_valid_b(array_6_io_d_out_0_valid_b),
    .io_d_out_1_a(array_6_io_d_out_1_a),
    .io_d_out_1_valid_a(array_6_io_d_out_1_valid_a),
    .io_d_out_1_b(array_6_io_d_out_1_b),
    .io_d_out_1_valid_b(array_6_io_d_out_1_valid_b),
    .io_d_out_2_a(array_6_io_d_out_2_a),
    .io_d_out_2_valid_a(array_6_io_d_out_2_valid_a),
    .io_d_out_2_b(array_6_io_d_out_2_b),
    .io_d_out_2_valid_b(array_6_io_d_out_2_valid_b),
    .io_d_out_3_a(array_6_io_d_out_3_a),
    .io_d_out_3_valid_a(array_6_io_d_out_3_valid_a),
    .io_d_out_3_b(array_6_io_d_out_3_b),
    .io_d_out_3_valid_b(array_6_io_d_out_3_valid_b),
    .io_d_out_4_a(array_6_io_d_out_4_a),
    .io_d_out_4_valid_a(array_6_io_d_out_4_valid_a),
    .io_d_out_4_b(array_6_io_d_out_4_b),
    .io_d_out_4_valid_b(array_6_io_d_out_4_valid_b),
    .io_d_out_5_a(array_6_io_d_out_5_a),
    .io_d_out_5_valid_a(array_6_io_d_out_5_valid_a),
    .io_d_out_5_b(array_6_io_d_out_5_b),
    .io_d_out_5_valid_b(array_6_io_d_out_5_valid_b),
    .io_d_out_6_a(array_6_io_d_out_6_a),
    .io_d_out_6_valid_a(array_6_io_d_out_6_valid_a),
    .io_d_out_6_b(array_6_io_d_out_6_b),
    .io_d_out_6_valid_b(array_6_io_d_out_6_valid_b),
    .io_d_out_7_a(array_6_io_d_out_7_a),
    .io_d_out_7_valid_a(array_6_io_d_out_7_valid_a),
    .io_d_out_7_b(array_6_io_d_out_7_b),
    .io_d_out_7_valid_b(array_6_io_d_out_7_valid_b),
    .io_d_out_8_a(array_6_io_d_out_8_a),
    .io_d_out_8_valid_a(array_6_io_d_out_8_valid_a),
    .io_d_out_8_b(array_6_io_d_out_8_b),
    .io_d_out_8_valid_b(array_6_io_d_out_8_valid_b),
    .io_d_out_9_a(array_6_io_d_out_9_a),
    .io_d_out_9_valid_a(array_6_io_d_out_9_valid_a),
    .io_d_out_9_b(array_6_io_d_out_9_b),
    .io_d_out_9_valid_b(array_6_io_d_out_9_valid_b),
    .io_d_out_10_a(array_6_io_d_out_10_a),
    .io_d_out_10_valid_a(array_6_io_d_out_10_valid_a),
    .io_d_out_10_b(array_6_io_d_out_10_b),
    .io_d_out_10_valid_b(array_6_io_d_out_10_valid_b),
    .io_d_out_11_a(array_6_io_d_out_11_a),
    .io_d_out_11_valid_a(array_6_io_d_out_11_valid_a),
    .io_d_out_11_b(array_6_io_d_out_11_b),
    .io_d_out_11_valid_b(array_6_io_d_out_11_valid_b),
    .io_d_out_12_a(array_6_io_d_out_12_a),
    .io_d_out_12_valid_a(array_6_io_d_out_12_valid_a),
    .io_d_out_12_b(array_6_io_d_out_12_b),
    .io_d_out_12_valid_b(array_6_io_d_out_12_valid_b),
    .io_d_out_13_a(array_6_io_d_out_13_a),
    .io_d_out_13_valid_a(array_6_io_d_out_13_valid_a),
    .io_d_out_13_b(array_6_io_d_out_13_b),
    .io_d_out_13_valid_b(array_6_io_d_out_13_valid_b),
    .io_d_out_14_a(array_6_io_d_out_14_a),
    .io_d_out_14_valid_a(array_6_io_d_out_14_valid_a),
    .io_d_out_14_b(array_6_io_d_out_14_b),
    .io_d_out_14_valid_b(array_6_io_d_out_14_valid_b),
    .io_d_out_15_a(array_6_io_d_out_15_a),
    .io_d_out_15_valid_a(array_6_io_d_out_15_valid_a),
    .io_d_out_15_b(array_6_io_d_out_15_b),
    .io_d_out_15_valid_b(array_6_io_d_out_15_valid_b),
    .io_d_out_16_a(array_6_io_d_out_16_a),
    .io_d_out_16_valid_a(array_6_io_d_out_16_valid_a),
    .io_d_out_16_b(array_6_io_d_out_16_b),
    .io_d_out_16_valid_b(array_6_io_d_out_16_valid_b),
    .io_d_out_17_a(array_6_io_d_out_17_a),
    .io_d_out_17_valid_a(array_6_io_d_out_17_valid_a),
    .io_d_out_17_b(array_6_io_d_out_17_b),
    .io_d_out_17_valid_b(array_6_io_d_out_17_valid_b),
    .io_d_out_18_a(array_6_io_d_out_18_a),
    .io_d_out_18_valid_a(array_6_io_d_out_18_valid_a),
    .io_d_out_18_b(array_6_io_d_out_18_b),
    .io_d_out_18_valid_b(array_6_io_d_out_18_valid_b),
    .io_d_out_19_a(array_6_io_d_out_19_a),
    .io_d_out_19_valid_a(array_6_io_d_out_19_valid_a),
    .io_d_out_19_b(array_6_io_d_out_19_b),
    .io_d_out_19_valid_b(array_6_io_d_out_19_valid_b),
    .io_d_out_20_a(array_6_io_d_out_20_a),
    .io_d_out_20_valid_a(array_6_io_d_out_20_valid_a),
    .io_d_out_20_b(array_6_io_d_out_20_b),
    .io_d_out_20_valid_b(array_6_io_d_out_20_valid_b),
    .io_d_out_21_a(array_6_io_d_out_21_a),
    .io_d_out_21_valid_a(array_6_io_d_out_21_valid_a),
    .io_d_out_21_b(array_6_io_d_out_21_b),
    .io_d_out_21_valid_b(array_6_io_d_out_21_valid_b),
    .io_d_out_22_a(array_6_io_d_out_22_a),
    .io_d_out_22_valid_a(array_6_io_d_out_22_valid_a),
    .io_d_out_22_b(array_6_io_d_out_22_b),
    .io_d_out_22_valid_b(array_6_io_d_out_22_valid_b),
    .io_d_out_23_a(array_6_io_d_out_23_a),
    .io_d_out_23_valid_a(array_6_io_d_out_23_valid_a),
    .io_d_out_23_b(array_6_io_d_out_23_b),
    .io_d_out_23_valid_b(array_6_io_d_out_23_valid_b),
    .io_d_out_24_a(array_6_io_d_out_24_a),
    .io_d_out_24_valid_a(array_6_io_d_out_24_valid_a),
    .io_d_out_24_b(array_6_io_d_out_24_b),
    .io_d_out_24_valid_b(array_6_io_d_out_24_valid_b),
    .io_d_out_25_a(array_6_io_d_out_25_a),
    .io_d_out_25_valid_a(array_6_io_d_out_25_valid_a),
    .io_d_out_25_b(array_6_io_d_out_25_b),
    .io_d_out_25_valid_b(array_6_io_d_out_25_valid_b),
    .io_d_out_26_a(array_6_io_d_out_26_a),
    .io_d_out_26_valid_a(array_6_io_d_out_26_valid_a),
    .io_d_out_26_b(array_6_io_d_out_26_b),
    .io_d_out_26_valid_b(array_6_io_d_out_26_valid_b),
    .io_d_out_27_a(array_6_io_d_out_27_a),
    .io_d_out_27_valid_a(array_6_io_d_out_27_valid_a),
    .io_d_out_27_b(array_6_io_d_out_27_b),
    .io_d_out_27_valid_b(array_6_io_d_out_27_valid_b),
    .io_d_out_28_a(array_6_io_d_out_28_a),
    .io_d_out_28_valid_a(array_6_io_d_out_28_valid_a),
    .io_d_out_28_b(array_6_io_d_out_28_b),
    .io_d_out_28_valid_b(array_6_io_d_out_28_valid_b),
    .io_d_out_29_a(array_6_io_d_out_29_a),
    .io_d_out_29_valid_a(array_6_io_d_out_29_valid_a),
    .io_d_out_29_b(array_6_io_d_out_29_b),
    .io_d_out_29_valid_b(array_6_io_d_out_29_valid_b),
    .io_d_out_30_a(array_6_io_d_out_30_a),
    .io_d_out_30_valid_a(array_6_io_d_out_30_valid_a),
    .io_d_out_30_b(array_6_io_d_out_30_b),
    .io_d_out_30_valid_b(array_6_io_d_out_30_valid_b),
    .io_d_out_31_a(array_6_io_d_out_31_a),
    .io_d_out_31_valid_a(array_6_io_d_out_31_valid_a),
    .io_d_out_31_b(array_6_io_d_out_31_b),
    .io_d_out_31_valid_b(array_6_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_6_io_wr_en_mem1),
    .io_wr_en_mem2(array_6_io_wr_en_mem2),
    .io_wr_en_mem3(array_6_io_wr_en_mem3),
    .io_wr_en_mem4(array_6_io_wr_en_mem4),
    .io_wr_en_mem5(array_6_io_wr_en_mem5),
    .io_wr_en_mem6(array_6_io_wr_en_mem6),
    .io_wr_instr_mem1(array_6_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_6_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_6_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_6_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_6_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_6_io_wr_instr_mem6),
    .io_PC1_in(array_6_io_PC1_in),
    .io_PC6_out(array_6_io_PC6_out),
    .io_Addr_in(array_6_io_Addr_in),
    .io_Addr_out(array_6_io_Addr_out)
  );
  BuildingBlockNew array_7 ( // @[BP.scala 45:51]
    .clock(array_7_clock),
    .reset(array_7_reset),
    .io_d_in_0_a(array_7_io_d_in_0_a),
    .io_d_in_0_valid_a(array_7_io_d_in_0_valid_a),
    .io_d_in_0_b(array_7_io_d_in_0_b),
    .io_d_in_0_valid_b(array_7_io_d_in_0_valid_b),
    .io_d_in_1_a(array_7_io_d_in_1_a),
    .io_d_in_1_valid_a(array_7_io_d_in_1_valid_a),
    .io_d_in_1_b(array_7_io_d_in_1_b),
    .io_d_in_1_valid_b(array_7_io_d_in_1_valid_b),
    .io_d_in_2_a(array_7_io_d_in_2_a),
    .io_d_in_2_valid_a(array_7_io_d_in_2_valid_a),
    .io_d_in_2_b(array_7_io_d_in_2_b),
    .io_d_in_2_valid_b(array_7_io_d_in_2_valid_b),
    .io_d_in_3_a(array_7_io_d_in_3_a),
    .io_d_in_3_valid_a(array_7_io_d_in_3_valid_a),
    .io_d_in_3_b(array_7_io_d_in_3_b),
    .io_d_in_3_valid_b(array_7_io_d_in_3_valid_b),
    .io_d_in_4_a(array_7_io_d_in_4_a),
    .io_d_in_4_valid_a(array_7_io_d_in_4_valid_a),
    .io_d_in_4_b(array_7_io_d_in_4_b),
    .io_d_in_4_valid_b(array_7_io_d_in_4_valid_b),
    .io_d_in_5_a(array_7_io_d_in_5_a),
    .io_d_in_5_valid_a(array_7_io_d_in_5_valid_a),
    .io_d_in_5_b(array_7_io_d_in_5_b),
    .io_d_in_5_valid_b(array_7_io_d_in_5_valid_b),
    .io_d_in_6_a(array_7_io_d_in_6_a),
    .io_d_in_6_valid_a(array_7_io_d_in_6_valid_a),
    .io_d_in_6_b(array_7_io_d_in_6_b),
    .io_d_in_6_valid_b(array_7_io_d_in_6_valid_b),
    .io_d_in_7_a(array_7_io_d_in_7_a),
    .io_d_in_7_valid_a(array_7_io_d_in_7_valid_a),
    .io_d_in_7_b(array_7_io_d_in_7_b),
    .io_d_in_7_valid_b(array_7_io_d_in_7_valid_b),
    .io_d_in_8_a(array_7_io_d_in_8_a),
    .io_d_in_8_valid_a(array_7_io_d_in_8_valid_a),
    .io_d_in_8_b(array_7_io_d_in_8_b),
    .io_d_in_8_valid_b(array_7_io_d_in_8_valid_b),
    .io_d_in_9_a(array_7_io_d_in_9_a),
    .io_d_in_9_valid_a(array_7_io_d_in_9_valid_a),
    .io_d_in_9_b(array_7_io_d_in_9_b),
    .io_d_in_9_valid_b(array_7_io_d_in_9_valid_b),
    .io_d_in_10_a(array_7_io_d_in_10_a),
    .io_d_in_10_valid_a(array_7_io_d_in_10_valid_a),
    .io_d_in_10_b(array_7_io_d_in_10_b),
    .io_d_in_10_valid_b(array_7_io_d_in_10_valid_b),
    .io_d_in_11_a(array_7_io_d_in_11_a),
    .io_d_in_11_valid_a(array_7_io_d_in_11_valid_a),
    .io_d_in_11_b(array_7_io_d_in_11_b),
    .io_d_in_11_valid_b(array_7_io_d_in_11_valid_b),
    .io_d_in_12_a(array_7_io_d_in_12_a),
    .io_d_in_12_valid_a(array_7_io_d_in_12_valid_a),
    .io_d_in_12_b(array_7_io_d_in_12_b),
    .io_d_in_12_valid_b(array_7_io_d_in_12_valid_b),
    .io_d_in_13_a(array_7_io_d_in_13_a),
    .io_d_in_13_valid_a(array_7_io_d_in_13_valid_a),
    .io_d_in_13_b(array_7_io_d_in_13_b),
    .io_d_in_13_valid_b(array_7_io_d_in_13_valid_b),
    .io_d_in_14_a(array_7_io_d_in_14_a),
    .io_d_in_14_valid_a(array_7_io_d_in_14_valid_a),
    .io_d_in_14_b(array_7_io_d_in_14_b),
    .io_d_in_14_valid_b(array_7_io_d_in_14_valid_b),
    .io_d_in_15_a(array_7_io_d_in_15_a),
    .io_d_in_15_valid_a(array_7_io_d_in_15_valid_a),
    .io_d_in_15_b(array_7_io_d_in_15_b),
    .io_d_in_15_valid_b(array_7_io_d_in_15_valid_b),
    .io_d_in_16_a(array_7_io_d_in_16_a),
    .io_d_in_16_valid_a(array_7_io_d_in_16_valid_a),
    .io_d_in_16_b(array_7_io_d_in_16_b),
    .io_d_in_16_valid_b(array_7_io_d_in_16_valid_b),
    .io_d_in_17_a(array_7_io_d_in_17_a),
    .io_d_in_17_valid_a(array_7_io_d_in_17_valid_a),
    .io_d_in_17_b(array_7_io_d_in_17_b),
    .io_d_in_17_valid_b(array_7_io_d_in_17_valid_b),
    .io_d_in_18_a(array_7_io_d_in_18_a),
    .io_d_in_18_valid_a(array_7_io_d_in_18_valid_a),
    .io_d_in_18_b(array_7_io_d_in_18_b),
    .io_d_in_18_valid_b(array_7_io_d_in_18_valid_b),
    .io_d_in_19_a(array_7_io_d_in_19_a),
    .io_d_in_19_valid_a(array_7_io_d_in_19_valid_a),
    .io_d_in_19_b(array_7_io_d_in_19_b),
    .io_d_in_19_valid_b(array_7_io_d_in_19_valid_b),
    .io_d_in_20_a(array_7_io_d_in_20_a),
    .io_d_in_20_valid_a(array_7_io_d_in_20_valid_a),
    .io_d_in_20_b(array_7_io_d_in_20_b),
    .io_d_in_20_valid_b(array_7_io_d_in_20_valid_b),
    .io_d_in_21_a(array_7_io_d_in_21_a),
    .io_d_in_21_valid_a(array_7_io_d_in_21_valid_a),
    .io_d_in_21_b(array_7_io_d_in_21_b),
    .io_d_in_21_valid_b(array_7_io_d_in_21_valid_b),
    .io_d_in_22_a(array_7_io_d_in_22_a),
    .io_d_in_22_valid_a(array_7_io_d_in_22_valid_a),
    .io_d_in_22_b(array_7_io_d_in_22_b),
    .io_d_in_22_valid_b(array_7_io_d_in_22_valid_b),
    .io_d_in_23_a(array_7_io_d_in_23_a),
    .io_d_in_23_valid_a(array_7_io_d_in_23_valid_a),
    .io_d_in_23_b(array_7_io_d_in_23_b),
    .io_d_in_23_valid_b(array_7_io_d_in_23_valid_b),
    .io_d_in_24_a(array_7_io_d_in_24_a),
    .io_d_in_24_valid_a(array_7_io_d_in_24_valid_a),
    .io_d_in_24_b(array_7_io_d_in_24_b),
    .io_d_in_24_valid_b(array_7_io_d_in_24_valid_b),
    .io_d_in_25_a(array_7_io_d_in_25_a),
    .io_d_in_25_valid_a(array_7_io_d_in_25_valid_a),
    .io_d_in_25_b(array_7_io_d_in_25_b),
    .io_d_in_25_valid_b(array_7_io_d_in_25_valid_b),
    .io_d_in_26_a(array_7_io_d_in_26_a),
    .io_d_in_26_valid_a(array_7_io_d_in_26_valid_a),
    .io_d_in_26_b(array_7_io_d_in_26_b),
    .io_d_in_26_valid_b(array_7_io_d_in_26_valid_b),
    .io_d_in_27_a(array_7_io_d_in_27_a),
    .io_d_in_27_valid_a(array_7_io_d_in_27_valid_a),
    .io_d_in_27_b(array_7_io_d_in_27_b),
    .io_d_in_27_valid_b(array_7_io_d_in_27_valid_b),
    .io_d_in_28_a(array_7_io_d_in_28_a),
    .io_d_in_28_valid_a(array_7_io_d_in_28_valid_a),
    .io_d_in_28_b(array_7_io_d_in_28_b),
    .io_d_in_28_valid_b(array_7_io_d_in_28_valid_b),
    .io_d_in_29_a(array_7_io_d_in_29_a),
    .io_d_in_29_valid_a(array_7_io_d_in_29_valid_a),
    .io_d_in_29_b(array_7_io_d_in_29_b),
    .io_d_in_29_valid_b(array_7_io_d_in_29_valid_b),
    .io_d_in_30_a(array_7_io_d_in_30_a),
    .io_d_in_30_valid_a(array_7_io_d_in_30_valid_a),
    .io_d_in_30_b(array_7_io_d_in_30_b),
    .io_d_in_30_valid_b(array_7_io_d_in_30_valid_b),
    .io_d_in_31_a(array_7_io_d_in_31_a),
    .io_d_in_31_valid_a(array_7_io_d_in_31_valid_a),
    .io_d_in_31_b(array_7_io_d_in_31_b),
    .io_d_in_31_valid_b(array_7_io_d_in_31_valid_b),
    .io_d_out_0_a(array_7_io_d_out_0_a),
    .io_d_out_0_valid_a(array_7_io_d_out_0_valid_a),
    .io_d_out_0_b(array_7_io_d_out_0_b),
    .io_d_out_0_valid_b(array_7_io_d_out_0_valid_b),
    .io_d_out_1_a(array_7_io_d_out_1_a),
    .io_d_out_1_valid_a(array_7_io_d_out_1_valid_a),
    .io_d_out_1_b(array_7_io_d_out_1_b),
    .io_d_out_1_valid_b(array_7_io_d_out_1_valid_b),
    .io_d_out_2_a(array_7_io_d_out_2_a),
    .io_d_out_2_valid_a(array_7_io_d_out_2_valid_a),
    .io_d_out_2_b(array_7_io_d_out_2_b),
    .io_d_out_2_valid_b(array_7_io_d_out_2_valid_b),
    .io_d_out_3_a(array_7_io_d_out_3_a),
    .io_d_out_3_valid_a(array_7_io_d_out_3_valid_a),
    .io_d_out_3_b(array_7_io_d_out_3_b),
    .io_d_out_3_valid_b(array_7_io_d_out_3_valid_b),
    .io_d_out_4_a(array_7_io_d_out_4_a),
    .io_d_out_4_valid_a(array_7_io_d_out_4_valid_a),
    .io_d_out_4_b(array_7_io_d_out_4_b),
    .io_d_out_4_valid_b(array_7_io_d_out_4_valid_b),
    .io_d_out_5_a(array_7_io_d_out_5_a),
    .io_d_out_5_valid_a(array_7_io_d_out_5_valid_a),
    .io_d_out_5_b(array_7_io_d_out_5_b),
    .io_d_out_5_valid_b(array_7_io_d_out_5_valid_b),
    .io_d_out_6_a(array_7_io_d_out_6_a),
    .io_d_out_6_valid_a(array_7_io_d_out_6_valid_a),
    .io_d_out_6_b(array_7_io_d_out_6_b),
    .io_d_out_6_valid_b(array_7_io_d_out_6_valid_b),
    .io_d_out_7_a(array_7_io_d_out_7_a),
    .io_d_out_7_valid_a(array_7_io_d_out_7_valid_a),
    .io_d_out_7_b(array_7_io_d_out_7_b),
    .io_d_out_7_valid_b(array_7_io_d_out_7_valid_b),
    .io_d_out_8_a(array_7_io_d_out_8_a),
    .io_d_out_8_valid_a(array_7_io_d_out_8_valid_a),
    .io_d_out_8_b(array_7_io_d_out_8_b),
    .io_d_out_8_valid_b(array_7_io_d_out_8_valid_b),
    .io_d_out_9_a(array_7_io_d_out_9_a),
    .io_d_out_9_valid_a(array_7_io_d_out_9_valid_a),
    .io_d_out_9_b(array_7_io_d_out_9_b),
    .io_d_out_9_valid_b(array_7_io_d_out_9_valid_b),
    .io_d_out_10_a(array_7_io_d_out_10_a),
    .io_d_out_10_valid_a(array_7_io_d_out_10_valid_a),
    .io_d_out_10_b(array_7_io_d_out_10_b),
    .io_d_out_10_valid_b(array_7_io_d_out_10_valid_b),
    .io_d_out_11_a(array_7_io_d_out_11_a),
    .io_d_out_11_valid_a(array_7_io_d_out_11_valid_a),
    .io_d_out_11_b(array_7_io_d_out_11_b),
    .io_d_out_11_valid_b(array_7_io_d_out_11_valid_b),
    .io_d_out_12_a(array_7_io_d_out_12_a),
    .io_d_out_12_valid_a(array_7_io_d_out_12_valid_a),
    .io_d_out_12_b(array_7_io_d_out_12_b),
    .io_d_out_12_valid_b(array_7_io_d_out_12_valid_b),
    .io_d_out_13_a(array_7_io_d_out_13_a),
    .io_d_out_13_valid_a(array_7_io_d_out_13_valid_a),
    .io_d_out_13_b(array_7_io_d_out_13_b),
    .io_d_out_13_valid_b(array_7_io_d_out_13_valid_b),
    .io_d_out_14_a(array_7_io_d_out_14_a),
    .io_d_out_14_valid_a(array_7_io_d_out_14_valid_a),
    .io_d_out_14_b(array_7_io_d_out_14_b),
    .io_d_out_14_valid_b(array_7_io_d_out_14_valid_b),
    .io_d_out_15_a(array_7_io_d_out_15_a),
    .io_d_out_15_valid_a(array_7_io_d_out_15_valid_a),
    .io_d_out_15_b(array_7_io_d_out_15_b),
    .io_d_out_15_valid_b(array_7_io_d_out_15_valid_b),
    .io_d_out_16_a(array_7_io_d_out_16_a),
    .io_d_out_16_valid_a(array_7_io_d_out_16_valid_a),
    .io_d_out_16_b(array_7_io_d_out_16_b),
    .io_d_out_16_valid_b(array_7_io_d_out_16_valid_b),
    .io_d_out_17_a(array_7_io_d_out_17_a),
    .io_d_out_17_valid_a(array_7_io_d_out_17_valid_a),
    .io_d_out_17_b(array_7_io_d_out_17_b),
    .io_d_out_17_valid_b(array_7_io_d_out_17_valid_b),
    .io_d_out_18_a(array_7_io_d_out_18_a),
    .io_d_out_18_valid_a(array_7_io_d_out_18_valid_a),
    .io_d_out_18_b(array_7_io_d_out_18_b),
    .io_d_out_18_valid_b(array_7_io_d_out_18_valid_b),
    .io_d_out_19_a(array_7_io_d_out_19_a),
    .io_d_out_19_valid_a(array_7_io_d_out_19_valid_a),
    .io_d_out_19_b(array_7_io_d_out_19_b),
    .io_d_out_19_valid_b(array_7_io_d_out_19_valid_b),
    .io_d_out_20_a(array_7_io_d_out_20_a),
    .io_d_out_20_valid_a(array_7_io_d_out_20_valid_a),
    .io_d_out_20_b(array_7_io_d_out_20_b),
    .io_d_out_20_valid_b(array_7_io_d_out_20_valid_b),
    .io_d_out_21_a(array_7_io_d_out_21_a),
    .io_d_out_21_valid_a(array_7_io_d_out_21_valid_a),
    .io_d_out_21_b(array_7_io_d_out_21_b),
    .io_d_out_21_valid_b(array_7_io_d_out_21_valid_b),
    .io_d_out_22_a(array_7_io_d_out_22_a),
    .io_d_out_22_valid_a(array_7_io_d_out_22_valid_a),
    .io_d_out_22_b(array_7_io_d_out_22_b),
    .io_d_out_22_valid_b(array_7_io_d_out_22_valid_b),
    .io_d_out_23_a(array_7_io_d_out_23_a),
    .io_d_out_23_valid_a(array_7_io_d_out_23_valid_a),
    .io_d_out_23_b(array_7_io_d_out_23_b),
    .io_d_out_23_valid_b(array_7_io_d_out_23_valid_b),
    .io_d_out_24_a(array_7_io_d_out_24_a),
    .io_d_out_24_valid_a(array_7_io_d_out_24_valid_a),
    .io_d_out_24_b(array_7_io_d_out_24_b),
    .io_d_out_24_valid_b(array_7_io_d_out_24_valid_b),
    .io_d_out_25_a(array_7_io_d_out_25_a),
    .io_d_out_25_valid_a(array_7_io_d_out_25_valid_a),
    .io_d_out_25_b(array_7_io_d_out_25_b),
    .io_d_out_25_valid_b(array_7_io_d_out_25_valid_b),
    .io_d_out_26_a(array_7_io_d_out_26_a),
    .io_d_out_26_valid_a(array_7_io_d_out_26_valid_a),
    .io_d_out_26_b(array_7_io_d_out_26_b),
    .io_d_out_26_valid_b(array_7_io_d_out_26_valid_b),
    .io_d_out_27_a(array_7_io_d_out_27_a),
    .io_d_out_27_valid_a(array_7_io_d_out_27_valid_a),
    .io_d_out_27_b(array_7_io_d_out_27_b),
    .io_d_out_27_valid_b(array_7_io_d_out_27_valid_b),
    .io_d_out_28_a(array_7_io_d_out_28_a),
    .io_d_out_28_valid_a(array_7_io_d_out_28_valid_a),
    .io_d_out_28_b(array_7_io_d_out_28_b),
    .io_d_out_28_valid_b(array_7_io_d_out_28_valid_b),
    .io_d_out_29_a(array_7_io_d_out_29_a),
    .io_d_out_29_valid_a(array_7_io_d_out_29_valid_a),
    .io_d_out_29_b(array_7_io_d_out_29_b),
    .io_d_out_29_valid_b(array_7_io_d_out_29_valid_b),
    .io_d_out_30_a(array_7_io_d_out_30_a),
    .io_d_out_30_valid_a(array_7_io_d_out_30_valid_a),
    .io_d_out_30_b(array_7_io_d_out_30_b),
    .io_d_out_30_valid_b(array_7_io_d_out_30_valid_b),
    .io_d_out_31_a(array_7_io_d_out_31_a),
    .io_d_out_31_valid_a(array_7_io_d_out_31_valid_a),
    .io_d_out_31_b(array_7_io_d_out_31_b),
    .io_d_out_31_valid_b(array_7_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_7_io_wr_en_mem1),
    .io_wr_en_mem2(array_7_io_wr_en_mem2),
    .io_wr_en_mem3(array_7_io_wr_en_mem3),
    .io_wr_en_mem4(array_7_io_wr_en_mem4),
    .io_wr_en_mem5(array_7_io_wr_en_mem5),
    .io_wr_en_mem6(array_7_io_wr_en_mem6),
    .io_wr_instr_mem1(array_7_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_7_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_7_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_7_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_7_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_7_io_wr_instr_mem6),
    .io_PC1_in(array_7_io_PC1_in),
    .io_PC6_out(array_7_io_PC6_out),
    .io_Addr_in(array_7_io_Addr_in),
    .io_Addr_out(array_7_io_Addr_out)
  );
  BuildingBlockNew array_8 ( // @[BP.scala 45:51]
    .clock(array_8_clock),
    .reset(array_8_reset),
    .io_d_in_0_a(array_8_io_d_in_0_a),
    .io_d_in_0_valid_a(array_8_io_d_in_0_valid_a),
    .io_d_in_0_b(array_8_io_d_in_0_b),
    .io_d_in_0_valid_b(array_8_io_d_in_0_valid_b),
    .io_d_in_1_a(array_8_io_d_in_1_a),
    .io_d_in_1_valid_a(array_8_io_d_in_1_valid_a),
    .io_d_in_1_b(array_8_io_d_in_1_b),
    .io_d_in_1_valid_b(array_8_io_d_in_1_valid_b),
    .io_d_in_2_a(array_8_io_d_in_2_a),
    .io_d_in_2_valid_a(array_8_io_d_in_2_valid_a),
    .io_d_in_2_b(array_8_io_d_in_2_b),
    .io_d_in_2_valid_b(array_8_io_d_in_2_valid_b),
    .io_d_in_3_a(array_8_io_d_in_3_a),
    .io_d_in_3_valid_a(array_8_io_d_in_3_valid_a),
    .io_d_in_3_b(array_8_io_d_in_3_b),
    .io_d_in_3_valid_b(array_8_io_d_in_3_valid_b),
    .io_d_in_4_a(array_8_io_d_in_4_a),
    .io_d_in_4_valid_a(array_8_io_d_in_4_valid_a),
    .io_d_in_4_b(array_8_io_d_in_4_b),
    .io_d_in_4_valid_b(array_8_io_d_in_4_valid_b),
    .io_d_in_5_a(array_8_io_d_in_5_a),
    .io_d_in_5_valid_a(array_8_io_d_in_5_valid_a),
    .io_d_in_5_b(array_8_io_d_in_5_b),
    .io_d_in_5_valid_b(array_8_io_d_in_5_valid_b),
    .io_d_in_6_a(array_8_io_d_in_6_a),
    .io_d_in_6_valid_a(array_8_io_d_in_6_valid_a),
    .io_d_in_6_b(array_8_io_d_in_6_b),
    .io_d_in_6_valid_b(array_8_io_d_in_6_valid_b),
    .io_d_in_7_a(array_8_io_d_in_7_a),
    .io_d_in_7_valid_a(array_8_io_d_in_7_valid_a),
    .io_d_in_7_b(array_8_io_d_in_7_b),
    .io_d_in_7_valid_b(array_8_io_d_in_7_valid_b),
    .io_d_in_8_a(array_8_io_d_in_8_a),
    .io_d_in_8_valid_a(array_8_io_d_in_8_valid_a),
    .io_d_in_8_b(array_8_io_d_in_8_b),
    .io_d_in_8_valid_b(array_8_io_d_in_8_valid_b),
    .io_d_in_9_a(array_8_io_d_in_9_a),
    .io_d_in_9_valid_a(array_8_io_d_in_9_valid_a),
    .io_d_in_9_b(array_8_io_d_in_9_b),
    .io_d_in_9_valid_b(array_8_io_d_in_9_valid_b),
    .io_d_in_10_a(array_8_io_d_in_10_a),
    .io_d_in_10_valid_a(array_8_io_d_in_10_valid_a),
    .io_d_in_10_b(array_8_io_d_in_10_b),
    .io_d_in_10_valid_b(array_8_io_d_in_10_valid_b),
    .io_d_in_11_a(array_8_io_d_in_11_a),
    .io_d_in_11_valid_a(array_8_io_d_in_11_valid_a),
    .io_d_in_11_b(array_8_io_d_in_11_b),
    .io_d_in_11_valid_b(array_8_io_d_in_11_valid_b),
    .io_d_in_12_a(array_8_io_d_in_12_a),
    .io_d_in_12_valid_a(array_8_io_d_in_12_valid_a),
    .io_d_in_12_b(array_8_io_d_in_12_b),
    .io_d_in_12_valid_b(array_8_io_d_in_12_valid_b),
    .io_d_in_13_a(array_8_io_d_in_13_a),
    .io_d_in_13_valid_a(array_8_io_d_in_13_valid_a),
    .io_d_in_13_b(array_8_io_d_in_13_b),
    .io_d_in_13_valid_b(array_8_io_d_in_13_valid_b),
    .io_d_in_14_a(array_8_io_d_in_14_a),
    .io_d_in_14_valid_a(array_8_io_d_in_14_valid_a),
    .io_d_in_14_b(array_8_io_d_in_14_b),
    .io_d_in_14_valid_b(array_8_io_d_in_14_valid_b),
    .io_d_in_15_a(array_8_io_d_in_15_a),
    .io_d_in_15_valid_a(array_8_io_d_in_15_valid_a),
    .io_d_in_15_b(array_8_io_d_in_15_b),
    .io_d_in_15_valid_b(array_8_io_d_in_15_valid_b),
    .io_d_in_16_a(array_8_io_d_in_16_a),
    .io_d_in_16_valid_a(array_8_io_d_in_16_valid_a),
    .io_d_in_16_b(array_8_io_d_in_16_b),
    .io_d_in_16_valid_b(array_8_io_d_in_16_valid_b),
    .io_d_in_17_a(array_8_io_d_in_17_a),
    .io_d_in_17_valid_a(array_8_io_d_in_17_valid_a),
    .io_d_in_17_b(array_8_io_d_in_17_b),
    .io_d_in_17_valid_b(array_8_io_d_in_17_valid_b),
    .io_d_in_18_a(array_8_io_d_in_18_a),
    .io_d_in_18_valid_a(array_8_io_d_in_18_valid_a),
    .io_d_in_18_b(array_8_io_d_in_18_b),
    .io_d_in_18_valid_b(array_8_io_d_in_18_valid_b),
    .io_d_in_19_a(array_8_io_d_in_19_a),
    .io_d_in_19_valid_a(array_8_io_d_in_19_valid_a),
    .io_d_in_19_b(array_8_io_d_in_19_b),
    .io_d_in_19_valid_b(array_8_io_d_in_19_valid_b),
    .io_d_in_20_a(array_8_io_d_in_20_a),
    .io_d_in_20_valid_a(array_8_io_d_in_20_valid_a),
    .io_d_in_20_b(array_8_io_d_in_20_b),
    .io_d_in_20_valid_b(array_8_io_d_in_20_valid_b),
    .io_d_in_21_a(array_8_io_d_in_21_a),
    .io_d_in_21_valid_a(array_8_io_d_in_21_valid_a),
    .io_d_in_21_b(array_8_io_d_in_21_b),
    .io_d_in_21_valid_b(array_8_io_d_in_21_valid_b),
    .io_d_in_22_a(array_8_io_d_in_22_a),
    .io_d_in_22_valid_a(array_8_io_d_in_22_valid_a),
    .io_d_in_22_b(array_8_io_d_in_22_b),
    .io_d_in_22_valid_b(array_8_io_d_in_22_valid_b),
    .io_d_in_23_a(array_8_io_d_in_23_a),
    .io_d_in_23_valid_a(array_8_io_d_in_23_valid_a),
    .io_d_in_23_b(array_8_io_d_in_23_b),
    .io_d_in_23_valid_b(array_8_io_d_in_23_valid_b),
    .io_d_in_24_a(array_8_io_d_in_24_a),
    .io_d_in_24_valid_a(array_8_io_d_in_24_valid_a),
    .io_d_in_24_b(array_8_io_d_in_24_b),
    .io_d_in_24_valid_b(array_8_io_d_in_24_valid_b),
    .io_d_in_25_a(array_8_io_d_in_25_a),
    .io_d_in_25_valid_a(array_8_io_d_in_25_valid_a),
    .io_d_in_25_b(array_8_io_d_in_25_b),
    .io_d_in_25_valid_b(array_8_io_d_in_25_valid_b),
    .io_d_in_26_a(array_8_io_d_in_26_a),
    .io_d_in_26_valid_a(array_8_io_d_in_26_valid_a),
    .io_d_in_26_b(array_8_io_d_in_26_b),
    .io_d_in_26_valid_b(array_8_io_d_in_26_valid_b),
    .io_d_in_27_a(array_8_io_d_in_27_a),
    .io_d_in_27_valid_a(array_8_io_d_in_27_valid_a),
    .io_d_in_27_b(array_8_io_d_in_27_b),
    .io_d_in_27_valid_b(array_8_io_d_in_27_valid_b),
    .io_d_in_28_a(array_8_io_d_in_28_a),
    .io_d_in_28_valid_a(array_8_io_d_in_28_valid_a),
    .io_d_in_28_b(array_8_io_d_in_28_b),
    .io_d_in_28_valid_b(array_8_io_d_in_28_valid_b),
    .io_d_in_29_a(array_8_io_d_in_29_a),
    .io_d_in_29_valid_a(array_8_io_d_in_29_valid_a),
    .io_d_in_29_b(array_8_io_d_in_29_b),
    .io_d_in_29_valid_b(array_8_io_d_in_29_valid_b),
    .io_d_in_30_a(array_8_io_d_in_30_a),
    .io_d_in_30_valid_a(array_8_io_d_in_30_valid_a),
    .io_d_in_30_b(array_8_io_d_in_30_b),
    .io_d_in_30_valid_b(array_8_io_d_in_30_valid_b),
    .io_d_in_31_a(array_8_io_d_in_31_a),
    .io_d_in_31_valid_a(array_8_io_d_in_31_valid_a),
    .io_d_in_31_b(array_8_io_d_in_31_b),
    .io_d_in_31_valid_b(array_8_io_d_in_31_valid_b),
    .io_d_out_0_a(array_8_io_d_out_0_a),
    .io_d_out_0_valid_a(array_8_io_d_out_0_valid_a),
    .io_d_out_0_b(array_8_io_d_out_0_b),
    .io_d_out_0_valid_b(array_8_io_d_out_0_valid_b),
    .io_d_out_1_a(array_8_io_d_out_1_a),
    .io_d_out_1_valid_a(array_8_io_d_out_1_valid_a),
    .io_d_out_1_b(array_8_io_d_out_1_b),
    .io_d_out_1_valid_b(array_8_io_d_out_1_valid_b),
    .io_d_out_2_a(array_8_io_d_out_2_a),
    .io_d_out_2_valid_a(array_8_io_d_out_2_valid_a),
    .io_d_out_2_b(array_8_io_d_out_2_b),
    .io_d_out_2_valid_b(array_8_io_d_out_2_valid_b),
    .io_d_out_3_a(array_8_io_d_out_3_a),
    .io_d_out_3_valid_a(array_8_io_d_out_3_valid_a),
    .io_d_out_3_b(array_8_io_d_out_3_b),
    .io_d_out_3_valid_b(array_8_io_d_out_3_valid_b),
    .io_d_out_4_a(array_8_io_d_out_4_a),
    .io_d_out_4_valid_a(array_8_io_d_out_4_valid_a),
    .io_d_out_4_b(array_8_io_d_out_4_b),
    .io_d_out_4_valid_b(array_8_io_d_out_4_valid_b),
    .io_d_out_5_a(array_8_io_d_out_5_a),
    .io_d_out_5_valid_a(array_8_io_d_out_5_valid_a),
    .io_d_out_5_b(array_8_io_d_out_5_b),
    .io_d_out_5_valid_b(array_8_io_d_out_5_valid_b),
    .io_d_out_6_a(array_8_io_d_out_6_a),
    .io_d_out_6_valid_a(array_8_io_d_out_6_valid_a),
    .io_d_out_6_b(array_8_io_d_out_6_b),
    .io_d_out_6_valid_b(array_8_io_d_out_6_valid_b),
    .io_d_out_7_a(array_8_io_d_out_7_a),
    .io_d_out_7_valid_a(array_8_io_d_out_7_valid_a),
    .io_d_out_7_b(array_8_io_d_out_7_b),
    .io_d_out_7_valid_b(array_8_io_d_out_7_valid_b),
    .io_d_out_8_a(array_8_io_d_out_8_a),
    .io_d_out_8_valid_a(array_8_io_d_out_8_valid_a),
    .io_d_out_8_b(array_8_io_d_out_8_b),
    .io_d_out_8_valid_b(array_8_io_d_out_8_valid_b),
    .io_d_out_9_a(array_8_io_d_out_9_a),
    .io_d_out_9_valid_a(array_8_io_d_out_9_valid_a),
    .io_d_out_9_b(array_8_io_d_out_9_b),
    .io_d_out_9_valid_b(array_8_io_d_out_9_valid_b),
    .io_d_out_10_a(array_8_io_d_out_10_a),
    .io_d_out_10_valid_a(array_8_io_d_out_10_valid_a),
    .io_d_out_10_b(array_8_io_d_out_10_b),
    .io_d_out_10_valid_b(array_8_io_d_out_10_valid_b),
    .io_d_out_11_a(array_8_io_d_out_11_a),
    .io_d_out_11_valid_a(array_8_io_d_out_11_valid_a),
    .io_d_out_11_b(array_8_io_d_out_11_b),
    .io_d_out_11_valid_b(array_8_io_d_out_11_valid_b),
    .io_d_out_12_a(array_8_io_d_out_12_a),
    .io_d_out_12_valid_a(array_8_io_d_out_12_valid_a),
    .io_d_out_12_b(array_8_io_d_out_12_b),
    .io_d_out_12_valid_b(array_8_io_d_out_12_valid_b),
    .io_d_out_13_a(array_8_io_d_out_13_a),
    .io_d_out_13_valid_a(array_8_io_d_out_13_valid_a),
    .io_d_out_13_b(array_8_io_d_out_13_b),
    .io_d_out_13_valid_b(array_8_io_d_out_13_valid_b),
    .io_d_out_14_a(array_8_io_d_out_14_a),
    .io_d_out_14_valid_a(array_8_io_d_out_14_valid_a),
    .io_d_out_14_b(array_8_io_d_out_14_b),
    .io_d_out_14_valid_b(array_8_io_d_out_14_valid_b),
    .io_d_out_15_a(array_8_io_d_out_15_a),
    .io_d_out_15_valid_a(array_8_io_d_out_15_valid_a),
    .io_d_out_15_b(array_8_io_d_out_15_b),
    .io_d_out_15_valid_b(array_8_io_d_out_15_valid_b),
    .io_d_out_16_a(array_8_io_d_out_16_a),
    .io_d_out_16_valid_a(array_8_io_d_out_16_valid_a),
    .io_d_out_16_b(array_8_io_d_out_16_b),
    .io_d_out_16_valid_b(array_8_io_d_out_16_valid_b),
    .io_d_out_17_a(array_8_io_d_out_17_a),
    .io_d_out_17_valid_a(array_8_io_d_out_17_valid_a),
    .io_d_out_17_b(array_8_io_d_out_17_b),
    .io_d_out_17_valid_b(array_8_io_d_out_17_valid_b),
    .io_d_out_18_a(array_8_io_d_out_18_a),
    .io_d_out_18_valid_a(array_8_io_d_out_18_valid_a),
    .io_d_out_18_b(array_8_io_d_out_18_b),
    .io_d_out_18_valid_b(array_8_io_d_out_18_valid_b),
    .io_d_out_19_a(array_8_io_d_out_19_a),
    .io_d_out_19_valid_a(array_8_io_d_out_19_valid_a),
    .io_d_out_19_b(array_8_io_d_out_19_b),
    .io_d_out_19_valid_b(array_8_io_d_out_19_valid_b),
    .io_d_out_20_a(array_8_io_d_out_20_a),
    .io_d_out_20_valid_a(array_8_io_d_out_20_valid_a),
    .io_d_out_20_b(array_8_io_d_out_20_b),
    .io_d_out_20_valid_b(array_8_io_d_out_20_valid_b),
    .io_d_out_21_a(array_8_io_d_out_21_a),
    .io_d_out_21_valid_a(array_8_io_d_out_21_valid_a),
    .io_d_out_21_b(array_8_io_d_out_21_b),
    .io_d_out_21_valid_b(array_8_io_d_out_21_valid_b),
    .io_d_out_22_a(array_8_io_d_out_22_a),
    .io_d_out_22_valid_a(array_8_io_d_out_22_valid_a),
    .io_d_out_22_b(array_8_io_d_out_22_b),
    .io_d_out_22_valid_b(array_8_io_d_out_22_valid_b),
    .io_d_out_23_a(array_8_io_d_out_23_a),
    .io_d_out_23_valid_a(array_8_io_d_out_23_valid_a),
    .io_d_out_23_b(array_8_io_d_out_23_b),
    .io_d_out_23_valid_b(array_8_io_d_out_23_valid_b),
    .io_d_out_24_a(array_8_io_d_out_24_a),
    .io_d_out_24_valid_a(array_8_io_d_out_24_valid_a),
    .io_d_out_24_b(array_8_io_d_out_24_b),
    .io_d_out_24_valid_b(array_8_io_d_out_24_valid_b),
    .io_d_out_25_a(array_8_io_d_out_25_a),
    .io_d_out_25_valid_a(array_8_io_d_out_25_valid_a),
    .io_d_out_25_b(array_8_io_d_out_25_b),
    .io_d_out_25_valid_b(array_8_io_d_out_25_valid_b),
    .io_d_out_26_a(array_8_io_d_out_26_a),
    .io_d_out_26_valid_a(array_8_io_d_out_26_valid_a),
    .io_d_out_26_b(array_8_io_d_out_26_b),
    .io_d_out_26_valid_b(array_8_io_d_out_26_valid_b),
    .io_d_out_27_a(array_8_io_d_out_27_a),
    .io_d_out_27_valid_a(array_8_io_d_out_27_valid_a),
    .io_d_out_27_b(array_8_io_d_out_27_b),
    .io_d_out_27_valid_b(array_8_io_d_out_27_valid_b),
    .io_d_out_28_a(array_8_io_d_out_28_a),
    .io_d_out_28_valid_a(array_8_io_d_out_28_valid_a),
    .io_d_out_28_b(array_8_io_d_out_28_b),
    .io_d_out_28_valid_b(array_8_io_d_out_28_valid_b),
    .io_d_out_29_a(array_8_io_d_out_29_a),
    .io_d_out_29_valid_a(array_8_io_d_out_29_valid_a),
    .io_d_out_29_b(array_8_io_d_out_29_b),
    .io_d_out_29_valid_b(array_8_io_d_out_29_valid_b),
    .io_d_out_30_a(array_8_io_d_out_30_a),
    .io_d_out_30_valid_a(array_8_io_d_out_30_valid_a),
    .io_d_out_30_b(array_8_io_d_out_30_b),
    .io_d_out_30_valid_b(array_8_io_d_out_30_valid_b),
    .io_d_out_31_a(array_8_io_d_out_31_a),
    .io_d_out_31_valid_a(array_8_io_d_out_31_valid_a),
    .io_d_out_31_b(array_8_io_d_out_31_b),
    .io_d_out_31_valid_b(array_8_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_8_io_wr_en_mem1),
    .io_wr_en_mem2(array_8_io_wr_en_mem2),
    .io_wr_en_mem3(array_8_io_wr_en_mem3),
    .io_wr_en_mem4(array_8_io_wr_en_mem4),
    .io_wr_en_mem5(array_8_io_wr_en_mem5),
    .io_wr_en_mem6(array_8_io_wr_en_mem6),
    .io_wr_instr_mem1(array_8_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_8_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_8_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_8_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_8_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_8_io_wr_instr_mem6),
    .io_PC1_in(array_8_io_PC1_in),
    .io_PC6_out(array_8_io_PC6_out),
    .io_Addr_in(array_8_io_Addr_in),
    .io_Addr_out(array_8_io_Addr_out)
  );
  BuildingBlockNew array_9 ( // @[BP.scala 45:51]
    .clock(array_9_clock),
    .reset(array_9_reset),
    .io_d_in_0_a(array_9_io_d_in_0_a),
    .io_d_in_0_valid_a(array_9_io_d_in_0_valid_a),
    .io_d_in_0_b(array_9_io_d_in_0_b),
    .io_d_in_0_valid_b(array_9_io_d_in_0_valid_b),
    .io_d_in_1_a(array_9_io_d_in_1_a),
    .io_d_in_1_valid_a(array_9_io_d_in_1_valid_a),
    .io_d_in_1_b(array_9_io_d_in_1_b),
    .io_d_in_1_valid_b(array_9_io_d_in_1_valid_b),
    .io_d_in_2_a(array_9_io_d_in_2_a),
    .io_d_in_2_valid_a(array_9_io_d_in_2_valid_a),
    .io_d_in_2_b(array_9_io_d_in_2_b),
    .io_d_in_2_valid_b(array_9_io_d_in_2_valid_b),
    .io_d_in_3_a(array_9_io_d_in_3_a),
    .io_d_in_3_valid_a(array_9_io_d_in_3_valid_a),
    .io_d_in_3_b(array_9_io_d_in_3_b),
    .io_d_in_3_valid_b(array_9_io_d_in_3_valid_b),
    .io_d_in_4_a(array_9_io_d_in_4_a),
    .io_d_in_4_valid_a(array_9_io_d_in_4_valid_a),
    .io_d_in_4_b(array_9_io_d_in_4_b),
    .io_d_in_4_valid_b(array_9_io_d_in_4_valid_b),
    .io_d_in_5_a(array_9_io_d_in_5_a),
    .io_d_in_5_valid_a(array_9_io_d_in_5_valid_a),
    .io_d_in_5_b(array_9_io_d_in_5_b),
    .io_d_in_5_valid_b(array_9_io_d_in_5_valid_b),
    .io_d_in_6_a(array_9_io_d_in_6_a),
    .io_d_in_6_valid_a(array_9_io_d_in_6_valid_a),
    .io_d_in_6_b(array_9_io_d_in_6_b),
    .io_d_in_6_valid_b(array_9_io_d_in_6_valid_b),
    .io_d_in_7_a(array_9_io_d_in_7_a),
    .io_d_in_7_valid_a(array_9_io_d_in_7_valid_a),
    .io_d_in_7_b(array_9_io_d_in_7_b),
    .io_d_in_7_valid_b(array_9_io_d_in_7_valid_b),
    .io_d_in_8_a(array_9_io_d_in_8_a),
    .io_d_in_8_valid_a(array_9_io_d_in_8_valid_a),
    .io_d_in_8_b(array_9_io_d_in_8_b),
    .io_d_in_8_valid_b(array_9_io_d_in_8_valid_b),
    .io_d_in_9_a(array_9_io_d_in_9_a),
    .io_d_in_9_valid_a(array_9_io_d_in_9_valid_a),
    .io_d_in_9_b(array_9_io_d_in_9_b),
    .io_d_in_9_valid_b(array_9_io_d_in_9_valid_b),
    .io_d_in_10_a(array_9_io_d_in_10_a),
    .io_d_in_10_valid_a(array_9_io_d_in_10_valid_a),
    .io_d_in_10_b(array_9_io_d_in_10_b),
    .io_d_in_10_valid_b(array_9_io_d_in_10_valid_b),
    .io_d_in_11_a(array_9_io_d_in_11_a),
    .io_d_in_11_valid_a(array_9_io_d_in_11_valid_a),
    .io_d_in_11_b(array_9_io_d_in_11_b),
    .io_d_in_11_valid_b(array_9_io_d_in_11_valid_b),
    .io_d_in_12_a(array_9_io_d_in_12_a),
    .io_d_in_12_valid_a(array_9_io_d_in_12_valid_a),
    .io_d_in_12_b(array_9_io_d_in_12_b),
    .io_d_in_12_valid_b(array_9_io_d_in_12_valid_b),
    .io_d_in_13_a(array_9_io_d_in_13_a),
    .io_d_in_13_valid_a(array_9_io_d_in_13_valid_a),
    .io_d_in_13_b(array_9_io_d_in_13_b),
    .io_d_in_13_valid_b(array_9_io_d_in_13_valid_b),
    .io_d_in_14_a(array_9_io_d_in_14_a),
    .io_d_in_14_valid_a(array_9_io_d_in_14_valid_a),
    .io_d_in_14_b(array_9_io_d_in_14_b),
    .io_d_in_14_valid_b(array_9_io_d_in_14_valid_b),
    .io_d_in_15_a(array_9_io_d_in_15_a),
    .io_d_in_15_valid_a(array_9_io_d_in_15_valid_a),
    .io_d_in_15_b(array_9_io_d_in_15_b),
    .io_d_in_15_valid_b(array_9_io_d_in_15_valid_b),
    .io_d_in_16_a(array_9_io_d_in_16_a),
    .io_d_in_16_valid_a(array_9_io_d_in_16_valid_a),
    .io_d_in_16_b(array_9_io_d_in_16_b),
    .io_d_in_16_valid_b(array_9_io_d_in_16_valid_b),
    .io_d_in_17_a(array_9_io_d_in_17_a),
    .io_d_in_17_valid_a(array_9_io_d_in_17_valid_a),
    .io_d_in_17_b(array_9_io_d_in_17_b),
    .io_d_in_17_valid_b(array_9_io_d_in_17_valid_b),
    .io_d_in_18_a(array_9_io_d_in_18_a),
    .io_d_in_18_valid_a(array_9_io_d_in_18_valid_a),
    .io_d_in_18_b(array_9_io_d_in_18_b),
    .io_d_in_18_valid_b(array_9_io_d_in_18_valid_b),
    .io_d_in_19_a(array_9_io_d_in_19_a),
    .io_d_in_19_valid_a(array_9_io_d_in_19_valid_a),
    .io_d_in_19_b(array_9_io_d_in_19_b),
    .io_d_in_19_valid_b(array_9_io_d_in_19_valid_b),
    .io_d_in_20_a(array_9_io_d_in_20_a),
    .io_d_in_20_valid_a(array_9_io_d_in_20_valid_a),
    .io_d_in_20_b(array_9_io_d_in_20_b),
    .io_d_in_20_valid_b(array_9_io_d_in_20_valid_b),
    .io_d_in_21_a(array_9_io_d_in_21_a),
    .io_d_in_21_valid_a(array_9_io_d_in_21_valid_a),
    .io_d_in_21_b(array_9_io_d_in_21_b),
    .io_d_in_21_valid_b(array_9_io_d_in_21_valid_b),
    .io_d_in_22_a(array_9_io_d_in_22_a),
    .io_d_in_22_valid_a(array_9_io_d_in_22_valid_a),
    .io_d_in_22_b(array_9_io_d_in_22_b),
    .io_d_in_22_valid_b(array_9_io_d_in_22_valid_b),
    .io_d_in_23_a(array_9_io_d_in_23_a),
    .io_d_in_23_valid_a(array_9_io_d_in_23_valid_a),
    .io_d_in_23_b(array_9_io_d_in_23_b),
    .io_d_in_23_valid_b(array_9_io_d_in_23_valid_b),
    .io_d_in_24_a(array_9_io_d_in_24_a),
    .io_d_in_24_valid_a(array_9_io_d_in_24_valid_a),
    .io_d_in_24_b(array_9_io_d_in_24_b),
    .io_d_in_24_valid_b(array_9_io_d_in_24_valid_b),
    .io_d_in_25_a(array_9_io_d_in_25_a),
    .io_d_in_25_valid_a(array_9_io_d_in_25_valid_a),
    .io_d_in_25_b(array_9_io_d_in_25_b),
    .io_d_in_25_valid_b(array_9_io_d_in_25_valid_b),
    .io_d_in_26_a(array_9_io_d_in_26_a),
    .io_d_in_26_valid_a(array_9_io_d_in_26_valid_a),
    .io_d_in_26_b(array_9_io_d_in_26_b),
    .io_d_in_26_valid_b(array_9_io_d_in_26_valid_b),
    .io_d_in_27_a(array_9_io_d_in_27_a),
    .io_d_in_27_valid_a(array_9_io_d_in_27_valid_a),
    .io_d_in_27_b(array_9_io_d_in_27_b),
    .io_d_in_27_valid_b(array_9_io_d_in_27_valid_b),
    .io_d_in_28_a(array_9_io_d_in_28_a),
    .io_d_in_28_valid_a(array_9_io_d_in_28_valid_a),
    .io_d_in_28_b(array_9_io_d_in_28_b),
    .io_d_in_28_valid_b(array_9_io_d_in_28_valid_b),
    .io_d_in_29_a(array_9_io_d_in_29_a),
    .io_d_in_29_valid_a(array_9_io_d_in_29_valid_a),
    .io_d_in_29_b(array_9_io_d_in_29_b),
    .io_d_in_29_valid_b(array_9_io_d_in_29_valid_b),
    .io_d_in_30_a(array_9_io_d_in_30_a),
    .io_d_in_30_valid_a(array_9_io_d_in_30_valid_a),
    .io_d_in_30_b(array_9_io_d_in_30_b),
    .io_d_in_30_valid_b(array_9_io_d_in_30_valid_b),
    .io_d_in_31_a(array_9_io_d_in_31_a),
    .io_d_in_31_valid_a(array_9_io_d_in_31_valid_a),
    .io_d_in_31_b(array_9_io_d_in_31_b),
    .io_d_in_31_valid_b(array_9_io_d_in_31_valid_b),
    .io_d_out_0_a(array_9_io_d_out_0_a),
    .io_d_out_0_valid_a(array_9_io_d_out_0_valid_a),
    .io_d_out_0_b(array_9_io_d_out_0_b),
    .io_d_out_0_valid_b(array_9_io_d_out_0_valid_b),
    .io_d_out_1_a(array_9_io_d_out_1_a),
    .io_d_out_1_valid_a(array_9_io_d_out_1_valid_a),
    .io_d_out_1_b(array_9_io_d_out_1_b),
    .io_d_out_1_valid_b(array_9_io_d_out_1_valid_b),
    .io_d_out_2_a(array_9_io_d_out_2_a),
    .io_d_out_2_valid_a(array_9_io_d_out_2_valid_a),
    .io_d_out_2_b(array_9_io_d_out_2_b),
    .io_d_out_2_valid_b(array_9_io_d_out_2_valid_b),
    .io_d_out_3_a(array_9_io_d_out_3_a),
    .io_d_out_3_valid_a(array_9_io_d_out_3_valid_a),
    .io_d_out_3_b(array_9_io_d_out_3_b),
    .io_d_out_3_valid_b(array_9_io_d_out_3_valid_b),
    .io_d_out_4_a(array_9_io_d_out_4_a),
    .io_d_out_4_valid_a(array_9_io_d_out_4_valid_a),
    .io_d_out_4_b(array_9_io_d_out_4_b),
    .io_d_out_4_valid_b(array_9_io_d_out_4_valid_b),
    .io_d_out_5_a(array_9_io_d_out_5_a),
    .io_d_out_5_valid_a(array_9_io_d_out_5_valid_a),
    .io_d_out_5_b(array_9_io_d_out_5_b),
    .io_d_out_5_valid_b(array_9_io_d_out_5_valid_b),
    .io_d_out_6_a(array_9_io_d_out_6_a),
    .io_d_out_6_valid_a(array_9_io_d_out_6_valid_a),
    .io_d_out_6_b(array_9_io_d_out_6_b),
    .io_d_out_6_valid_b(array_9_io_d_out_6_valid_b),
    .io_d_out_7_a(array_9_io_d_out_7_a),
    .io_d_out_7_valid_a(array_9_io_d_out_7_valid_a),
    .io_d_out_7_b(array_9_io_d_out_7_b),
    .io_d_out_7_valid_b(array_9_io_d_out_7_valid_b),
    .io_d_out_8_a(array_9_io_d_out_8_a),
    .io_d_out_8_valid_a(array_9_io_d_out_8_valid_a),
    .io_d_out_8_b(array_9_io_d_out_8_b),
    .io_d_out_8_valid_b(array_9_io_d_out_8_valid_b),
    .io_d_out_9_a(array_9_io_d_out_9_a),
    .io_d_out_9_valid_a(array_9_io_d_out_9_valid_a),
    .io_d_out_9_b(array_9_io_d_out_9_b),
    .io_d_out_9_valid_b(array_9_io_d_out_9_valid_b),
    .io_d_out_10_a(array_9_io_d_out_10_a),
    .io_d_out_10_valid_a(array_9_io_d_out_10_valid_a),
    .io_d_out_10_b(array_9_io_d_out_10_b),
    .io_d_out_10_valid_b(array_9_io_d_out_10_valid_b),
    .io_d_out_11_a(array_9_io_d_out_11_a),
    .io_d_out_11_valid_a(array_9_io_d_out_11_valid_a),
    .io_d_out_11_b(array_9_io_d_out_11_b),
    .io_d_out_11_valid_b(array_9_io_d_out_11_valid_b),
    .io_d_out_12_a(array_9_io_d_out_12_a),
    .io_d_out_12_valid_a(array_9_io_d_out_12_valid_a),
    .io_d_out_12_b(array_9_io_d_out_12_b),
    .io_d_out_12_valid_b(array_9_io_d_out_12_valid_b),
    .io_d_out_13_a(array_9_io_d_out_13_a),
    .io_d_out_13_valid_a(array_9_io_d_out_13_valid_a),
    .io_d_out_13_b(array_9_io_d_out_13_b),
    .io_d_out_13_valid_b(array_9_io_d_out_13_valid_b),
    .io_d_out_14_a(array_9_io_d_out_14_a),
    .io_d_out_14_valid_a(array_9_io_d_out_14_valid_a),
    .io_d_out_14_b(array_9_io_d_out_14_b),
    .io_d_out_14_valid_b(array_9_io_d_out_14_valid_b),
    .io_d_out_15_a(array_9_io_d_out_15_a),
    .io_d_out_15_valid_a(array_9_io_d_out_15_valid_a),
    .io_d_out_15_b(array_9_io_d_out_15_b),
    .io_d_out_15_valid_b(array_9_io_d_out_15_valid_b),
    .io_d_out_16_a(array_9_io_d_out_16_a),
    .io_d_out_16_valid_a(array_9_io_d_out_16_valid_a),
    .io_d_out_16_b(array_9_io_d_out_16_b),
    .io_d_out_16_valid_b(array_9_io_d_out_16_valid_b),
    .io_d_out_17_a(array_9_io_d_out_17_a),
    .io_d_out_17_valid_a(array_9_io_d_out_17_valid_a),
    .io_d_out_17_b(array_9_io_d_out_17_b),
    .io_d_out_17_valid_b(array_9_io_d_out_17_valid_b),
    .io_d_out_18_a(array_9_io_d_out_18_a),
    .io_d_out_18_valid_a(array_9_io_d_out_18_valid_a),
    .io_d_out_18_b(array_9_io_d_out_18_b),
    .io_d_out_18_valid_b(array_9_io_d_out_18_valid_b),
    .io_d_out_19_a(array_9_io_d_out_19_a),
    .io_d_out_19_valid_a(array_9_io_d_out_19_valid_a),
    .io_d_out_19_b(array_9_io_d_out_19_b),
    .io_d_out_19_valid_b(array_9_io_d_out_19_valid_b),
    .io_d_out_20_a(array_9_io_d_out_20_a),
    .io_d_out_20_valid_a(array_9_io_d_out_20_valid_a),
    .io_d_out_20_b(array_9_io_d_out_20_b),
    .io_d_out_20_valid_b(array_9_io_d_out_20_valid_b),
    .io_d_out_21_a(array_9_io_d_out_21_a),
    .io_d_out_21_valid_a(array_9_io_d_out_21_valid_a),
    .io_d_out_21_b(array_9_io_d_out_21_b),
    .io_d_out_21_valid_b(array_9_io_d_out_21_valid_b),
    .io_d_out_22_a(array_9_io_d_out_22_a),
    .io_d_out_22_valid_a(array_9_io_d_out_22_valid_a),
    .io_d_out_22_b(array_9_io_d_out_22_b),
    .io_d_out_22_valid_b(array_9_io_d_out_22_valid_b),
    .io_d_out_23_a(array_9_io_d_out_23_a),
    .io_d_out_23_valid_a(array_9_io_d_out_23_valid_a),
    .io_d_out_23_b(array_9_io_d_out_23_b),
    .io_d_out_23_valid_b(array_9_io_d_out_23_valid_b),
    .io_d_out_24_a(array_9_io_d_out_24_a),
    .io_d_out_24_valid_a(array_9_io_d_out_24_valid_a),
    .io_d_out_24_b(array_9_io_d_out_24_b),
    .io_d_out_24_valid_b(array_9_io_d_out_24_valid_b),
    .io_d_out_25_a(array_9_io_d_out_25_a),
    .io_d_out_25_valid_a(array_9_io_d_out_25_valid_a),
    .io_d_out_25_b(array_9_io_d_out_25_b),
    .io_d_out_25_valid_b(array_9_io_d_out_25_valid_b),
    .io_d_out_26_a(array_9_io_d_out_26_a),
    .io_d_out_26_valid_a(array_9_io_d_out_26_valid_a),
    .io_d_out_26_b(array_9_io_d_out_26_b),
    .io_d_out_26_valid_b(array_9_io_d_out_26_valid_b),
    .io_d_out_27_a(array_9_io_d_out_27_a),
    .io_d_out_27_valid_a(array_9_io_d_out_27_valid_a),
    .io_d_out_27_b(array_9_io_d_out_27_b),
    .io_d_out_27_valid_b(array_9_io_d_out_27_valid_b),
    .io_d_out_28_a(array_9_io_d_out_28_a),
    .io_d_out_28_valid_a(array_9_io_d_out_28_valid_a),
    .io_d_out_28_b(array_9_io_d_out_28_b),
    .io_d_out_28_valid_b(array_9_io_d_out_28_valid_b),
    .io_d_out_29_a(array_9_io_d_out_29_a),
    .io_d_out_29_valid_a(array_9_io_d_out_29_valid_a),
    .io_d_out_29_b(array_9_io_d_out_29_b),
    .io_d_out_29_valid_b(array_9_io_d_out_29_valid_b),
    .io_d_out_30_a(array_9_io_d_out_30_a),
    .io_d_out_30_valid_a(array_9_io_d_out_30_valid_a),
    .io_d_out_30_b(array_9_io_d_out_30_b),
    .io_d_out_30_valid_b(array_9_io_d_out_30_valid_b),
    .io_d_out_31_a(array_9_io_d_out_31_a),
    .io_d_out_31_valid_a(array_9_io_d_out_31_valid_a),
    .io_d_out_31_b(array_9_io_d_out_31_b),
    .io_d_out_31_valid_b(array_9_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_9_io_wr_en_mem1),
    .io_wr_en_mem2(array_9_io_wr_en_mem2),
    .io_wr_en_mem3(array_9_io_wr_en_mem3),
    .io_wr_en_mem4(array_9_io_wr_en_mem4),
    .io_wr_en_mem5(array_9_io_wr_en_mem5),
    .io_wr_en_mem6(array_9_io_wr_en_mem6),
    .io_wr_instr_mem1(array_9_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_9_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_9_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_9_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_9_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_9_io_wr_instr_mem6),
    .io_PC1_in(array_9_io_PC1_in),
    .io_PC6_out(array_9_io_PC6_out),
    .io_Addr_in(array_9_io_Addr_in),
    .io_Addr_out(array_9_io_Addr_out)
  );
  BuildingBlockNew array_10 ( // @[BP.scala 45:51]
    .clock(array_10_clock),
    .reset(array_10_reset),
    .io_d_in_0_a(array_10_io_d_in_0_a),
    .io_d_in_0_valid_a(array_10_io_d_in_0_valid_a),
    .io_d_in_0_b(array_10_io_d_in_0_b),
    .io_d_in_0_valid_b(array_10_io_d_in_0_valid_b),
    .io_d_in_1_a(array_10_io_d_in_1_a),
    .io_d_in_1_valid_a(array_10_io_d_in_1_valid_a),
    .io_d_in_1_b(array_10_io_d_in_1_b),
    .io_d_in_1_valid_b(array_10_io_d_in_1_valid_b),
    .io_d_in_2_a(array_10_io_d_in_2_a),
    .io_d_in_2_valid_a(array_10_io_d_in_2_valid_a),
    .io_d_in_2_b(array_10_io_d_in_2_b),
    .io_d_in_2_valid_b(array_10_io_d_in_2_valid_b),
    .io_d_in_3_a(array_10_io_d_in_3_a),
    .io_d_in_3_valid_a(array_10_io_d_in_3_valid_a),
    .io_d_in_3_b(array_10_io_d_in_3_b),
    .io_d_in_3_valid_b(array_10_io_d_in_3_valid_b),
    .io_d_in_4_a(array_10_io_d_in_4_a),
    .io_d_in_4_valid_a(array_10_io_d_in_4_valid_a),
    .io_d_in_4_b(array_10_io_d_in_4_b),
    .io_d_in_4_valid_b(array_10_io_d_in_4_valid_b),
    .io_d_in_5_a(array_10_io_d_in_5_a),
    .io_d_in_5_valid_a(array_10_io_d_in_5_valid_a),
    .io_d_in_5_b(array_10_io_d_in_5_b),
    .io_d_in_5_valid_b(array_10_io_d_in_5_valid_b),
    .io_d_in_6_a(array_10_io_d_in_6_a),
    .io_d_in_6_valid_a(array_10_io_d_in_6_valid_a),
    .io_d_in_6_b(array_10_io_d_in_6_b),
    .io_d_in_6_valid_b(array_10_io_d_in_6_valid_b),
    .io_d_in_7_a(array_10_io_d_in_7_a),
    .io_d_in_7_valid_a(array_10_io_d_in_7_valid_a),
    .io_d_in_7_b(array_10_io_d_in_7_b),
    .io_d_in_7_valid_b(array_10_io_d_in_7_valid_b),
    .io_d_in_8_a(array_10_io_d_in_8_a),
    .io_d_in_8_valid_a(array_10_io_d_in_8_valid_a),
    .io_d_in_8_b(array_10_io_d_in_8_b),
    .io_d_in_8_valid_b(array_10_io_d_in_8_valid_b),
    .io_d_in_9_a(array_10_io_d_in_9_a),
    .io_d_in_9_valid_a(array_10_io_d_in_9_valid_a),
    .io_d_in_9_b(array_10_io_d_in_9_b),
    .io_d_in_9_valid_b(array_10_io_d_in_9_valid_b),
    .io_d_in_10_a(array_10_io_d_in_10_a),
    .io_d_in_10_valid_a(array_10_io_d_in_10_valid_a),
    .io_d_in_10_b(array_10_io_d_in_10_b),
    .io_d_in_10_valid_b(array_10_io_d_in_10_valid_b),
    .io_d_in_11_a(array_10_io_d_in_11_a),
    .io_d_in_11_valid_a(array_10_io_d_in_11_valid_a),
    .io_d_in_11_b(array_10_io_d_in_11_b),
    .io_d_in_11_valid_b(array_10_io_d_in_11_valid_b),
    .io_d_in_12_a(array_10_io_d_in_12_a),
    .io_d_in_12_valid_a(array_10_io_d_in_12_valid_a),
    .io_d_in_12_b(array_10_io_d_in_12_b),
    .io_d_in_12_valid_b(array_10_io_d_in_12_valid_b),
    .io_d_in_13_a(array_10_io_d_in_13_a),
    .io_d_in_13_valid_a(array_10_io_d_in_13_valid_a),
    .io_d_in_13_b(array_10_io_d_in_13_b),
    .io_d_in_13_valid_b(array_10_io_d_in_13_valid_b),
    .io_d_in_14_a(array_10_io_d_in_14_a),
    .io_d_in_14_valid_a(array_10_io_d_in_14_valid_a),
    .io_d_in_14_b(array_10_io_d_in_14_b),
    .io_d_in_14_valid_b(array_10_io_d_in_14_valid_b),
    .io_d_in_15_a(array_10_io_d_in_15_a),
    .io_d_in_15_valid_a(array_10_io_d_in_15_valid_a),
    .io_d_in_15_b(array_10_io_d_in_15_b),
    .io_d_in_15_valid_b(array_10_io_d_in_15_valid_b),
    .io_d_in_16_a(array_10_io_d_in_16_a),
    .io_d_in_16_valid_a(array_10_io_d_in_16_valid_a),
    .io_d_in_16_b(array_10_io_d_in_16_b),
    .io_d_in_16_valid_b(array_10_io_d_in_16_valid_b),
    .io_d_in_17_a(array_10_io_d_in_17_a),
    .io_d_in_17_valid_a(array_10_io_d_in_17_valid_a),
    .io_d_in_17_b(array_10_io_d_in_17_b),
    .io_d_in_17_valid_b(array_10_io_d_in_17_valid_b),
    .io_d_in_18_a(array_10_io_d_in_18_a),
    .io_d_in_18_valid_a(array_10_io_d_in_18_valid_a),
    .io_d_in_18_b(array_10_io_d_in_18_b),
    .io_d_in_18_valid_b(array_10_io_d_in_18_valid_b),
    .io_d_in_19_a(array_10_io_d_in_19_a),
    .io_d_in_19_valid_a(array_10_io_d_in_19_valid_a),
    .io_d_in_19_b(array_10_io_d_in_19_b),
    .io_d_in_19_valid_b(array_10_io_d_in_19_valid_b),
    .io_d_in_20_a(array_10_io_d_in_20_a),
    .io_d_in_20_valid_a(array_10_io_d_in_20_valid_a),
    .io_d_in_20_b(array_10_io_d_in_20_b),
    .io_d_in_20_valid_b(array_10_io_d_in_20_valid_b),
    .io_d_in_21_a(array_10_io_d_in_21_a),
    .io_d_in_21_valid_a(array_10_io_d_in_21_valid_a),
    .io_d_in_21_b(array_10_io_d_in_21_b),
    .io_d_in_21_valid_b(array_10_io_d_in_21_valid_b),
    .io_d_in_22_a(array_10_io_d_in_22_a),
    .io_d_in_22_valid_a(array_10_io_d_in_22_valid_a),
    .io_d_in_22_b(array_10_io_d_in_22_b),
    .io_d_in_22_valid_b(array_10_io_d_in_22_valid_b),
    .io_d_in_23_a(array_10_io_d_in_23_a),
    .io_d_in_23_valid_a(array_10_io_d_in_23_valid_a),
    .io_d_in_23_b(array_10_io_d_in_23_b),
    .io_d_in_23_valid_b(array_10_io_d_in_23_valid_b),
    .io_d_in_24_a(array_10_io_d_in_24_a),
    .io_d_in_24_valid_a(array_10_io_d_in_24_valid_a),
    .io_d_in_24_b(array_10_io_d_in_24_b),
    .io_d_in_24_valid_b(array_10_io_d_in_24_valid_b),
    .io_d_in_25_a(array_10_io_d_in_25_a),
    .io_d_in_25_valid_a(array_10_io_d_in_25_valid_a),
    .io_d_in_25_b(array_10_io_d_in_25_b),
    .io_d_in_25_valid_b(array_10_io_d_in_25_valid_b),
    .io_d_in_26_a(array_10_io_d_in_26_a),
    .io_d_in_26_valid_a(array_10_io_d_in_26_valid_a),
    .io_d_in_26_b(array_10_io_d_in_26_b),
    .io_d_in_26_valid_b(array_10_io_d_in_26_valid_b),
    .io_d_in_27_a(array_10_io_d_in_27_a),
    .io_d_in_27_valid_a(array_10_io_d_in_27_valid_a),
    .io_d_in_27_b(array_10_io_d_in_27_b),
    .io_d_in_27_valid_b(array_10_io_d_in_27_valid_b),
    .io_d_in_28_a(array_10_io_d_in_28_a),
    .io_d_in_28_valid_a(array_10_io_d_in_28_valid_a),
    .io_d_in_28_b(array_10_io_d_in_28_b),
    .io_d_in_28_valid_b(array_10_io_d_in_28_valid_b),
    .io_d_in_29_a(array_10_io_d_in_29_a),
    .io_d_in_29_valid_a(array_10_io_d_in_29_valid_a),
    .io_d_in_29_b(array_10_io_d_in_29_b),
    .io_d_in_29_valid_b(array_10_io_d_in_29_valid_b),
    .io_d_in_30_a(array_10_io_d_in_30_a),
    .io_d_in_30_valid_a(array_10_io_d_in_30_valid_a),
    .io_d_in_30_b(array_10_io_d_in_30_b),
    .io_d_in_30_valid_b(array_10_io_d_in_30_valid_b),
    .io_d_in_31_a(array_10_io_d_in_31_a),
    .io_d_in_31_valid_a(array_10_io_d_in_31_valid_a),
    .io_d_in_31_b(array_10_io_d_in_31_b),
    .io_d_in_31_valid_b(array_10_io_d_in_31_valid_b),
    .io_d_out_0_a(array_10_io_d_out_0_a),
    .io_d_out_0_valid_a(array_10_io_d_out_0_valid_a),
    .io_d_out_0_b(array_10_io_d_out_0_b),
    .io_d_out_0_valid_b(array_10_io_d_out_0_valid_b),
    .io_d_out_1_a(array_10_io_d_out_1_a),
    .io_d_out_1_valid_a(array_10_io_d_out_1_valid_a),
    .io_d_out_1_b(array_10_io_d_out_1_b),
    .io_d_out_1_valid_b(array_10_io_d_out_1_valid_b),
    .io_d_out_2_a(array_10_io_d_out_2_a),
    .io_d_out_2_valid_a(array_10_io_d_out_2_valid_a),
    .io_d_out_2_b(array_10_io_d_out_2_b),
    .io_d_out_2_valid_b(array_10_io_d_out_2_valid_b),
    .io_d_out_3_a(array_10_io_d_out_3_a),
    .io_d_out_3_valid_a(array_10_io_d_out_3_valid_a),
    .io_d_out_3_b(array_10_io_d_out_3_b),
    .io_d_out_3_valid_b(array_10_io_d_out_3_valid_b),
    .io_d_out_4_a(array_10_io_d_out_4_a),
    .io_d_out_4_valid_a(array_10_io_d_out_4_valid_a),
    .io_d_out_4_b(array_10_io_d_out_4_b),
    .io_d_out_4_valid_b(array_10_io_d_out_4_valid_b),
    .io_d_out_5_a(array_10_io_d_out_5_a),
    .io_d_out_5_valid_a(array_10_io_d_out_5_valid_a),
    .io_d_out_5_b(array_10_io_d_out_5_b),
    .io_d_out_5_valid_b(array_10_io_d_out_5_valid_b),
    .io_d_out_6_a(array_10_io_d_out_6_a),
    .io_d_out_6_valid_a(array_10_io_d_out_6_valid_a),
    .io_d_out_6_b(array_10_io_d_out_6_b),
    .io_d_out_6_valid_b(array_10_io_d_out_6_valid_b),
    .io_d_out_7_a(array_10_io_d_out_7_a),
    .io_d_out_7_valid_a(array_10_io_d_out_7_valid_a),
    .io_d_out_7_b(array_10_io_d_out_7_b),
    .io_d_out_7_valid_b(array_10_io_d_out_7_valid_b),
    .io_d_out_8_a(array_10_io_d_out_8_a),
    .io_d_out_8_valid_a(array_10_io_d_out_8_valid_a),
    .io_d_out_8_b(array_10_io_d_out_8_b),
    .io_d_out_8_valid_b(array_10_io_d_out_8_valid_b),
    .io_d_out_9_a(array_10_io_d_out_9_a),
    .io_d_out_9_valid_a(array_10_io_d_out_9_valid_a),
    .io_d_out_9_b(array_10_io_d_out_9_b),
    .io_d_out_9_valid_b(array_10_io_d_out_9_valid_b),
    .io_d_out_10_a(array_10_io_d_out_10_a),
    .io_d_out_10_valid_a(array_10_io_d_out_10_valid_a),
    .io_d_out_10_b(array_10_io_d_out_10_b),
    .io_d_out_10_valid_b(array_10_io_d_out_10_valid_b),
    .io_d_out_11_a(array_10_io_d_out_11_a),
    .io_d_out_11_valid_a(array_10_io_d_out_11_valid_a),
    .io_d_out_11_b(array_10_io_d_out_11_b),
    .io_d_out_11_valid_b(array_10_io_d_out_11_valid_b),
    .io_d_out_12_a(array_10_io_d_out_12_a),
    .io_d_out_12_valid_a(array_10_io_d_out_12_valid_a),
    .io_d_out_12_b(array_10_io_d_out_12_b),
    .io_d_out_12_valid_b(array_10_io_d_out_12_valid_b),
    .io_d_out_13_a(array_10_io_d_out_13_a),
    .io_d_out_13_valid_a(array_10_io_d_out_13_valid_a),
    .io_d_out_13_b(array_10_io_d_out_13_b),
    .io_d_out_13_valid_b(array_10_io_d_out_13_valid_b),
    .io_d_out_14_a(array_10_io_d_out_14_a),
    .io_d_out_14_valid_a(array_10_io_d_out_14_valid_a),
    .io_d_out_14_b(array_10_io_d_out_14_b),
    .io_d_out_14_valid_b(array_10_io_d_out_14_valid_b),
    .io_d_out_15_a(array_10_io_d_out_15_a),
    .io_d_out_15_valid_a(array_10_io_d_out_15_valid_a),
    .io_d_out_15_b(array_10_io_d_out_15_b),
    .io_d_out_15_valid_b(array_10_io_d_out_15_valid_b),
    .io_d_out_16_a(array_10_io_d_out_16_a),
    .io_d_out_16_valid_a(array_10_io_d_out_16_valid_a),
    .io_d_out_16_b(array_10_io_d_out_16_b),
    .io_d_out_16_valid_b(array_10_io_d_out_16_valid_b),
    .io_d_out_17_a(array_10_io_d_out_17_a),
    .io_d_out_17_valid_a(array_10_io_d_out_17_valid_a),
    .io_d_out_17_b(array_10_io_d_out_17_b),
    .io_d_out_17_valid_b(array_10_io_d_out_17_valid_b),
    .io_d_out_18_a(array_10_io_d_out_18_a),
    .io_d_out_18_valid_a(array_10_io_d_out_18_valid_a),
    .io_d_out_18_b(array_10_io_d_out_18_b),
    .io_d_out_18_valid_b(array_10_io_d_out_18_valid_b),
    .io_d_out_19_a(array_10_io_d_out_19_a),
    .io_d_out_19_valid_a(array_10_io_d_out_19_valid_a),
    .io_d_out_19_b(array_10_io_d_out_19_b),
    .io_d_out_19_valid_b(array_10_io_d_out_19_valid_b),
    .io_d_out_20_a(array_10_io_d_out_20_a),
    .io_d_out_20_valid_a(array_10_io_d_out_20_valid_a),
    .io_d_out_20_b(array_10_io_d_out_20_b),
    .io_d_out_20_valid_b(array_10_io_d_out_20_valid_b),
    .io_d_out_21_a(array_10_io_d_out_21_a),
    .io_d_out_21_valid_a(array_10_io_d_out_21_valid_a),
    .io_d_out_21_b(array_10_io_d_out_21_b),
    .io_d_out_21_valid_b(array_10_io_d_out_21_valid_b),
    .io_d_out_22_a(array_10_io_d_out_22_a),
    .io_d_out_22_valid_a(array_10_io_d_out_22_valid_a),
    .io_d_out_22_b(array_10_io_d_out_22_b),
    .io_d_out_22_valid_b(array_10_io_d_out_22_valid_b),
    .io_d_out_23_a(array_10_io_d_out_23_a),
    .io_d_out_23_valid_a(array_10_io_d_out_23_valid_a),
    .io_d_out_23_b(array_10_io_d_out_23_b),
    .io_d_out_23_valid_b(array_10_io_d_out_23_valid_b),
    .io_d_out_24_a(array_10_io_d_out_24_a),
    .io_d_out_24_valid_a(array_10_io_d_out_24_valid_a),
    .io_d_out_24_b(array_10_io_d_out_24_b),
    .io_d_out_24_valid_b(array_10_io_d_out_24_valid_b),
    .io_d_out_25_a(array_10_io_d_out_25_a),
    .io_d_out_25_valid_a(array_10_io_d_out_25_valid_a),
    .io_d_out_25_b(array_10_io_d_out_25_b),
    .io_d_out_25_valid_b(array_10_io_d_out_25_valid_b),
    .io_d_out_26_a(array_10_io_d_out_26_a),
    .io_d_out_26_valid_a(array_10_io_d_out_26_valid_a),
    .io_d_out_26_b(array_10_io_d_out_26_b),
    .io_d_out_26_valid_b(array_10_io_d_out_26_valid_b),
    .io_d_out_27_a(array_10_io_d_out_27_a),
    .io_d_out_27_valid_a(array_10_io_d_out_27_valid_a),
    .io_d_out_27_b(array_10_io_d_out_27_b),
    .io_d_out_27_valid_b(array_10_io_d_out_27_valid_b),
    .io_d_out_28_a(array_10_io_d_out_28_a),
    .io_d_out_28_valid_a(array_10_io_d_out_28_valid_a),
    .io_d_out_28_b(array_10_io_d_out_28_b),
    .io_d_out_28_valid_b(array_10_io_d_out_28_valid_b),
    .io_d_out_29_a(array_10_io_d_out_29_a),
    .io_d_out_29_valid_a(array_10_io_d_out_29_valid_a),
    .io_d_out_29_b(array_10_io_d_out_29_b),
    .io_d_out_29_valid_b(array_10_io_d_out_29_valid_b),
    .io_d_out_30_a(array_10_io_d_out_30_a),
    .io_d_out_30_valid_a(array_10_io_d_out_30_valid_a),
    .io_d_out_30_b(array_10_io_d_out_30_b),
    .io_d_out_30_valid_b(array_10_io_d_out_30_valid_b),
    .io_d_out_31_a(array_10_io_d_out_31_a),
    .io_d_out_31_valid_a(array_10_io_d_out_31_valid_a),
    .io_d_out_31_b(array_10_io_d_out_31_b),
    .io_d_out_31_valid_b(array_10_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_10_io_wr_en_mem1),
    .io_wr_en_mem2(array_10_io_wr_en_mem2),
    .io_wr_en_mem3(array_10_io_wr_en_mem3),
    .io_wr_en_mem4(array_10_io_wr_en_mem4),
    .io_wr_en_mem5(array_10_io_wr_en_mem5),
    .io_wr_en_mem6(array_10_io_wr_en_mem6),
    .io_wr_instr_mem1(array_10_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_10_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_10_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_10_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_10_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_10_io_wr_instr_mem6),
    .io_PC1_in(array_10_io_PC1_in),
    .io_PC6_out(array_10_io_PC6_out),
    .io_Addr_in(array_10_io_Addr_in),
    .io_Addr_out(array_10_io_Addr_out)
  );
  BuildingBlockNew array_11 ( // @[BP.scala 45:51]
    .clock(array_11_clock),
    .reset(array_11_reset),
    .io_d_in_0_a(array_11_io_d_in_0_a),
    .io_d_in_0_valid_a(array_11_io_d_in_0_valid_a),
    .io_d_in_0_b(array_11_io_d_in_0_b),
    .io_d_in_0_valid_b(array_11_io_d_in_0_valid_b),
    .io_d_in_1_a(array_11_io_d_in_1_a),
    .io_d_in_1_valid_a(array_11_io_d_in_1_valid_a),
    .io_d_in_1_b(array_11_io_d_in_1_b),
    .io_d_in_1_valid_b(array_11_io_d_in_1_valid_b),
    .io_d_in_2_a(array_11_io_d_in_2_a),
    .io_d_in_2_valid_a(array_11_io_d_in_2_valid_a),
    .io_d_in_2_b(array_11_io_d_in_2_b),
    .io_d_in_2_valid_b(array_11_io_d_in_2_valid_b),
    .io_d_in_3_a(array_11_io_d_in_3_a),
    .io_d_in_3_valid_a(array_11_io_d_in_3_valid_a),
    .io_d_in_3_b(array_11_io_d_in_3_b),
    .io_d_in_3_valid_b(array_11_io_d_in_3_valid_b),
    .io_d_in_4_a(array_11_io_d_in_4_a),
    .io_d_in_4_valid_a(array_11_io_d_in_4_valid_a),
    .io_d_in_4_b(array_11_io_d_in_4_b),
    .io_d_in_4_valid_b(array_11_io_d_in_4_valid_b),
    .io_d_in_5_a(array_11_io_d_in_5_a),
    .io_d_in_5_valid_a(array_11_io_d_in_5_valid_a),
    .io_d_in_5_b(array_11_io_d_in_5_b),
    .io_d_in_5_valid_b(array_11_io_d_in_5_valid_b),
    .io_d_in_6_a(array_11_io_d_in_6_a),
    .io_d_in_6_valid_a(array_11_io_d_in_6_valid_a),
    .io_d_in_6_b(array_11_io_d_in_6_b),
    .io_d_in_6_valid_b(array_11_io_d_in_6_valid_b),
    .io_d_in_7_a(array_11_io_d_in_7_a),
    .io_d_in_7_valid_a(array_11_io_d_in_7_valid_a),
    .io_d_in_7_b(array_11_io_d_in_7_b),
    .io_d_in_7_valid_b(array_11_io_d_in_7_valid_b),
    .io_d_in_8_a(array_11_io_d_in_8_a),
    .io_d_in_8_valid_a(array_11_io_d_in_8_valid_a),
    .io_d_in_8_b(array_11_io_d_in_8_b),
    .io_d_in_8_valid_b(array_11_io_d_in_8_valid_b),
    .io_d_in_9_a(array_11_io_d_in_9_a),
    .io_d_in_9_valid_a(array_11_io_d_in_9_valid_a),
    .io_d_in_9_b(array_11_io_d_in_9_b),
    .io_d_in_9_valid_b(array_11_io_d_in_9_valid_b),
    .io_d_in_10_a(array_11_io_d_in_10_a),
    .io_d_in_10_valid_a(array_11_io_d_in_10_valid_a),
    .io_d_in_10_b(array_11_io_d_in_10_b),
    .io_d_in_10_valid_b(array_11_io_d_in_10_valid_b),
    .io_d_in_11_a(array_11_io_d_in_11_a),
    .io_d_in_11_valid_a(array_11_io_d_in_11_valid_a),
    .io_d_in_11_b(array_11_io_d_in_11_b),
    .io_d_in_11_valid_b(array_11_io_d_in_11_valid_b),
    .io_d_in_12_a(array_11_io_d_in_12_a),
    .io_d_in_12_valid_a(array_11_io_d_in_12_valid_a),
    .io_d_in_12_b(array_11_io_d_in_12_b),
    .io_d_in_12_valid_b(array_11_io_d_in_12_valid_b),
    .io_d_in_13_a(array_11_io_d_in_13_a),
    .io_d_in_13_valid_a(array_11_io_d_in_13_valid_a),
    .io_d_in_13_b(array_11_io_d_in_13_b),
    .io_d_in_13_valid_b(array_11_io_d_in_13_valid_b),
    .io_d_in_14_a(array_11_io_d_in_14_a),
    .io_d_in_14_valid_a(array_11_io_d_in_14_valid_a),
    .io_d_in_14_b(array_11_io_d_in_14_b),
    .io_d_in_14_valid_b(array_11_io_d_in_14_valid_b),
    .io_d_in_15_a(array_11_io_d_in_15_a),
    .io_d_in_15_valid_a(array_11_io_d_in_15_valid_a),
    .io_d_in_15_b(array_11_io_d_in_15_b),
    .io_d_in_15_valid_b(array_11_io_d_in_15_valid_b),
    .io_d_in_16_a(array_11_io_d_in_16_a),
    .io_d_in_16_valid_a(array_11_io_d_in_16_valid_a),
    .io_d_in_16_b(array_11_io_d_in_16_b),
    .io_d_in_16_valid_b(array_11_io_d_in_16_valid_b),
    .io_d_in_17_a(array_11_io_d_in_17_a),
    .io_d_in_17_valid_a(array_11_io_d_in_17_valid_a),
    .io_d_in_17_b(array_11_io_d_in_17_b),
    .io_d_in_17_valid_b(array_11_io_d_in_17_valid_b),
    .io_d_in_18_a(array_11_io_d_in_18_a),
    .io_d_in_18_valid_a(array_11_io_d_in_18_valid_a),
    .io_d_in_18_b(array_11_io_d_in_18_b),
    .io_d_in_18_valid_b(array_11_io_d_in_18_valid_b),
    .io_d_in_19_a(array_11_io_d_in_19_a),
    .io_d_in_19_valid_a(array_11_io_d_in_19_valid_a),
    .io_d_in_19_b(array_11_io_d_in_19_b),
    .io_d_in_19_valid_b(array_11_io_d_in_19_valid_b),
    .io_d_in_20_a(array_11_io_d_in_20_a),
    .io_d_in_20_valid_a(array_11_io_d_in_20_valid_a),
    .io_d_in_20_b(array_11_io_d_in_20_b),
    .io_d_in_20_valid_b(array_11_io_d_in_20_valid_b),
    .io_d_in_21_a(array_11_io_d_in_21_a),
    .io_d_in_21_valid_a(array_11_io_d_in_21_valid_a),
    .io_d_in_21_b(array_11_io_d_in_21_b),
    .io_d_in_21_valid_b(array_11_io_d_in_21_valid_b),
    .io_d_in_22_a(array_11_io_d_in_22_a),
    .io_d_in_22_valid_a(array_11_io_d_in_22_valid_a),
    .io_d_in_22_b(array_11_io_d_in_22_b),
    .io_d_in_22_valid_b(array_11_io_d_in_22_valid_b),
    .io_d_in_23_a(array_11_io_d_in_23_a),
    .io_d_in_23_valid_a(array_11_io_d_in_23_valid_a),
    .io_d_in_23_b(array_11_io_d_in_23_b),
    .io_d_in_23_valid_b(array_11_io_d_in_23_valid_b),
    .io_d_in_24_a(array_11_io_d_in_24_a),
    .io_d_in_24_valid_a(array_11_io_d_in_24_valid_a),
    .io_d_in_24_b(array_11_io_d_in_24_b),
    .io_d_in_24_valid_b(array_11_io_d_in_24_valid_b),
    .io_d_in_25_a(array_11_io_d_in_25_a),
    .io_d_in_25_valid_a(array_11_io_d_in_25_valid_a),
    .io_d_in_25_b(array_11_io_d_in_25_b),
    .io_d_in_25_valid_b(array_11_io_d_in_25_valid_b),
    .io_d_in_26_a(array_11_io_d_in_26_a),
    .io_d_in_26_valid_a(array_11_io_d_in_26_valid_a),
    .io_d_in_26_b(array_11_io_d_in_26_b),
    .io_d_in_26_valid_b(array_11_io_d_in_26_valid_b),
    .io_d_in_27_a(array_11_io_d_in_27_a),
    .io_d_in_27_valid_a(array_11_io_d_in_27_valid_a),
    .io_d_in_27_b(array_11_io_d_in_27_b),
    .io_d_in_27_valid_b(array_11_io_d_in_27_valid_b),
    .io_d_in_28_a(array_11_io_d_in_28_a),
    .io_d_in_28_valid_a(array_11_io_d_in_28_valid_a),
    .io_d_in_28_b(array_11_io_d_in_28_b),
    .io_d_in_28_valid_b(array_11_io_d_in_28_valid_b),
    .io_d_in_29_a(array_11_io_d_in_29_a),
    .io_d_in_29_valid_a(array_11_io_d_in_29_valid_a),
    .io_d_in_29_b(array_11_io_d_in_29_b),
    .io_d_in_29_valid_b(array_11_io_d_in_29_valid_b),
    .io_d_in_30_a(array_11_io_d_in_30_a),
    .io_d_in_30_valid_a(array_11_io_d_in_30_valid_a),
    .io_d_in_30_b(array_11_io_d_in_30_b),
    .io_d_in_30_valid_b(array_11_io_d_in_30_valid_b),
    .io_d_in_31_a(array_11_io_d_in_31_a),
    .io_d_in_31_valid_a(array_11_io_d_in_31_valid_a),
    .io_d_in_31_b(array_11_io_d_in_31_b),
    .io_d_in_31_valid_b(array_11_io_d_in_31_valid_b),
    .io_d_out_0_a(array_11_io_d_out_0_a),
    .io_d_out_0_valid_a(array_11_io_d_out_0_valid_a),
    .io_d_out_0_b(array_11_io_d_out_0_b),
    .io_d_out_0_valid_b(array_11_io_d_out_0_valid_b),
    .io_d_out_1_a(array_11_io_d_out_1_a),
    .io_d_out_1_valid_a(array_11_io_d_out_1_valid_a),
    .io_d_out_1_b(array_11_io_d_out_1_b),
    .io_d_out_1_valid_b(array_11_io_d_out_1_valid_b),
    .io_d_out_2_a(array_11_io_d_out_2_a),
    .io_d_out_2_valid_a(array_11_io_d_out_2_valid_a),
    .io_d_out_2_b(array_11_io_d_out_2_b),
    .io_d_out_2_valid_b(array_11_io_d_out_2_valid_b),
    .io_d_out_3_a(array_11_io_d_out_3_a),
    .io_d_out_3_valid_a(array_11_io_d_out_3_valid_a),
    .io_d_out_3_b(array_11_io_d_out_3_b),
    .io_d_out_3_valid_b(array_11_io_d_out_3_valid_b),
    .io_d_out_4_a(array_11_io_d_out_4_a),
    .io_d_out_4_valid_a(array_11_io_d_out_4_valid_a),
    .io_d_out_4_b(array_11_io_d_out_4_b),
    .io_d_out_4_valid_b(array_11_io_d_out_4_valid_b),
    .io_d_out_5_a(array_11_io_d_out_5_a),
    .io_d_out_5_valid_a(array_11_io_d_out_5_valid_a),
    .io_d_out_5_b(array_11_io_d_out_5_b),
    .io_d_out_5_valid_b(array_11_io_d_out_5_valid_b),
    .io_d_out_6_a(array_11_io_d_out_6_a),
    .io_d_out_6_valid_a(array_11_io_d_out_6_valid_a),
    .io_d_out_6_b(array_11_io_d_out_6_b),
    .io_d_out_6_valid_b(array_11_io_d_out_6_valid_b),
    .io_d_out_7_a(array_11_io_d_out_7_a),
    .io_d_out_7_valid_a(array_11_io_d_out_7_valid_a),
    .io_d_out_7_b(array_11_io_d_out_7_b),
    .io_d_out_7_valid_b(array_11_io_d_out_7_valid_b),
    .io_d_out_8_a(array_11_io_d_out_8_a),
    .io_d_out_8_valid_a(array_11_io_d_out_8_valid_a),
    .io_d_out_8_b(array_11_io_d_out_8_b),
    .io_d_out_8_valid_b(array_11_io_d_out_8_valid_b),
    .io_d_out_9_a(array_11_io_d_out_9_a),
    .io_d_out_9_valid_a(array_11_io_d_out_9_valid_a),
    .io_d_out_9_b(array_11_io_d_out_9_b),
    .io_d_out_9_valid_b(array_11_io_d_out_9_valid_b),
    .io_d_out_10_a(array_11_io_d_out_10_a),
    .io_d_out_10_valid_a(array_11_io_d_out_10_valid_a),
    .io_d_out_10_b(array_11_io_d_out_10_b),
    .io_d_out_10_valid_b(array_11_io_d_out_10_valid_b),
    .io_d_out_11_a(array_11_io_d_out_11_a),
    .io_d_out_11_valid_a(array_11_io_d_out_11_valid_a),
    .io_d_out_11_b(array_11_io_d_out_11_b),
    .io_d_out_11_valid_b(array_11_io_d_out_11_valid_b),
    .io_d_out_12_a(array_11_io_d_out_12_a),
    .io_d_out_12_valid_a(array_11_io_d_out_12_valid_a),
    .io_d_out_12_b(array_11_io_d_out_12_b),
    .io_d_out_12_valid_b(array_11_io_d_out_12_valid_b),
    .io_d_out_13_a(array_11_io_d_out_13_a),
    .io_d_out_13_valid_a(array_11_io_d_out_13_valid_a),
    .io_d_out_13_b(array_11_io_d_out_13_b),
    .io_d_out_13_valid_b(array_11_io_d_out_13_valid_b),
    .io_d_out_14_a(array_11_io_d_out_14_a),
    .io_d_out_14_valid_a(array_11_io_d_out_14_valid_a),
    .io_d_out_14_b(array_11_io_d_out_14_b),
    .io_d_out_14_valid_b(array_11_io_d_out_14_valid_b),
    .io_d_out_15_a(array_11_io_d_out_15_a),
    .io_d_out_15_valid_a(array_11_io_d_out_15_valid_a),
    .io_d_out_15_b(array_11_io_d_out_15_b),
    .io_d_out_15_valid_b(array_11_io_d_out_15_valid_b),
    .io_d_out_16_a(array_11_io_d_out_16_a),
    .io_d_out_16_valid_a(array_11_io_d_out_16_valid_a),
    .io_d_out_16_b(array_11_io_d_out_16_b),
    .io_d_out_16_valid_b(array_11_io_d_out_16_valid_b),
    .io_d_out_17_a(array_11_io_d_out_17_a),
    .io_d_out_17_valid_a(array_11_io_d_out_17_valid_a),
    .io_d_out_17_b(array_11_io_d_out_17_b),
    .io_d_out_17_valid_b(array_11_io_d_out_17_valid_b),
    .io_d_out_18_a(array_11_io_d_out_18_a),
    .io_d_out_18_valid_a(array_11_io_d_out_18_valid_a),
    .io_d_out_18_b(array_11_io_d_out_18_b),
    .io_d_out_18_valid_b(array_11_io_d_out_18_valid_b),
    .io_d_out_19_a(array_11_io_d_out_19_a),
    .io_d_out_19_valid_a(array_11_io_d_out_19_valid_a),
    .io_d_out_19_b(array_11_io_d_out_19_b),
    .io_d_out_19_valid_b(array_11_io_d_out_19_valid_b),
    .io_d_out_20_a(array_11_io_d_out_20_a),
    .io_d_out_20_valid_a(array_11_io_d_out_20_valid_a),
    .io_d_out_20_b(array_11_io_d_out_20_b),
    .io_d_out_20_valid_b(array_11_io_d_out_20_valid_b),
    .io_d_out_21_a(array_11_io_d_out_21_a),
    .io_d_out_21_valid_a(array_11_io_d_out_21_valid_a),
    .io_d_out_21_b(array_11_io_d_out_21_b),
    .io_d_out_21_valid_b(array_11_io_d_out_21_valid_b),
    .io_d_out_22_a(array_11_io_d_out_22_a),
    .io_d_out_22_valid_a(array_11_io_d_out_22_valid_a),
    .io_d_out_22_b(array_11_io_d_out_22_b),
    .io_d_out_22_valid_b(array_11_io_d_out_22_valid_b),
    .io_d_out_23_a(array_11_io_d_out_23_a),
    .io_d_out_23_valid_a(array_11_io_d_out_23_valid_a),
    .io_d_out_23_b(array_11_io_d_out_23_b),
    .io_d_out_23_valid_b(array_11_io_d_out_23_valid_b),
    .io_d_out_24_a(array_11_io_d_out_24_a),
    .io_d_out_24_valid_a(array_11_io_d_out_24_valid_a),
    .io_d_out_24_b(array_11_io_d_out_24_b),
    .io_d_out_24_valid_b(array_11_io_d_out_24_valid_b),
    .io_d_out_25_a(array_11_io_d_out_25_a),
    .io_d_out_25_valid_a(array_11_io_d_out_25_valid_a),
    .io_d_out_25_b(array_11_io_d_out_25_b),
    .io_d_out_25_valid_b(array_11_io_d_out_25_valid_b),
    .io_d_out_26_a(array_11_io_d_out_26_a),
    .io_d_out_26_valid_a(array_11_io_d_out_26_valid_a),
    .io_d_out_26_b(array_11_io_d_out_26_b),
    .io_d_out_26_valid_b(array_11_io_d_out_26_valid_b),
    .io_d_out_27_a(array_11_io_d_out_27_a),
    .io_d_out_27_valid_a(array_11_io_d_out_27_valid_a),
    .io_d_out_27_b(array_11_io_d_out_27_b),
    .io_d_out_27_valid_b(array_11_io_d_out_27_valid_b),
    .io_d_out_28_a(array_11_io_d_out_28_a),
    .io_d_out_28_valid_a(array_11_io_d_out_28_valid_a),
    .io_d_out_28_b(array_11_io_d_out_28_b),
    .io_d_out_28_valid_b(array_11_io_d_out_28_valid_b),
    .io_d_out_29_a(array_11_io_d_out_29_a),
    .io_d_out_29_valid_a(array_11_io_d_out_29_valid_a),
    .io_d_out_29_b(array_11_io_d_out_29_b),
    .io_d_out_29_valid_b(array_11_io_d_out_29_valid_b),
    .io_d_out_30_a(array_11_io_d_out_30_a),
    .io_d_out_30_valid_a(array_11_io_d_out_30_valid_a),
    .io_d_out_30_b(array_11_io_d_out_30_b),
    .io_d_out_30_valid_b(array_11_io_d_out_30_valid_b),
    .io_d_out_31_a(array_11_io_d_out_31_a),
    .io_d_out_31_valid_a(array_11_io_d_out_31_valid_a),
    .io_d_out_31_b(array_11_io_d_out_31_b),
    .io_d_out_31_valid_b(array_11_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_11_io_wr_en_mem1),
    .io_wr_en_mem2(array_11_io_wr_en_mem2),
    .io_wr_en_mem3(array_11_io_wr_en_mem3),
    .io_wr_en_mem4(array_11_io_wr_en_mem4),
    .io_wr_en_mem5(array_11_io_wr_en_mem5),
    .io_wr_en_mem6(array_11_io_wr_en_mem6),
    .io_wr_instr_mem1(array_11_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_11_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_11_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_11_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_11_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_11_io_wr_instr_mem6),
    .io_PC1_in(array_11_io_PC1_in),
    .io_PC6_out(array_11_io_PC6_out),
    .io_Addr_in(array_11_io_Addr_in),
    .io_Addr_out(array_11_io_Addr_out)
  );
  BuildingBlockNew array_12 ( // @[BP.scala 45:51]
    .clock(array_12_clock),
    .reset(array_12_reset),
    .io_d_in_0_a(array_12_io_d_in_0_a),
    .io_d_in_0_valid_a(array_12_io_d_in_0_valid_a),
    .io_d_in_0_b(array_12_io_d_in_0_b),
    .io_d_in_0_valid_b(array_12_io_d_in_0_valid_b),
    .io_d_in_1_a(array_12_io_d_in_1_a),
    .io_d_in_1_valid_a(array_12_io_d_in_1_valid_a),
    .io_d_in_1_b(array_12_io_d_in_1_b),
    .io_d_in_1_valid_b(array_12_io_d_in_1_valid_b),
    .io_d_in_2_a(array_12_io_d_in_2_a),
    .io_d_in_2_valid_a(array_12_io_d_in_2_valid_a),
    .io_d_in_2_b(array_12_io_d_in_2_b),
    .io_d_in_2_valid_b(array_12_io_d_in_2_valid_b),
    .io_d_in_3_a(array_12_io_d_in_3_a),
    .io_d_in_3_valid_a(array_12_io_d_in_3_valid_a),
    .io_d_in_3_b(array_12_io_d_in_3_b),
    .io_d_in_3_valid_b(array_12_io_d_in_3_valid_b),
    .io_d_in_4_a(array_12_io_d_in_4_a),
    .io_d_in_4_valid_a(array_12_io_d_in_4_valid_a),
    .io_d_in_4_b(array_12_io_d_in_4_b),
    .io_d_in_4_valid_b(array_12_io_d_in_4_valid_b),
    .io_d_in_5_a(array_12_io_d_in_5_a),
    .io_d_in_5_valid_a(array_12_io_d_in_5_valid_a),
    .io_d_in_5_b(array_12_io_d_in_5_b),
    .io_d_in_5_valid_b(array_12_io_d_in_5_valid_b),
    .io_d_in_6_a(array_12_io_d_in_6_a),
    .io_d_in_6_valid_a(array_12_io_d_in_6_valid_a),
    .io_d_in_6_b(array_12_io_d_in_6_b),
    .io_d_in_6_valid_b(array_12_io_d_in_6_valid_b),
    .io_d_in_7_a(array_12_io_d_in_7_a),
    .io_d_in_7_valid_a(array_12_io_d_in_7_valid_a),
    .io_d_in_7_b(array_12_io_d_in_7_b),
    .io_d_in_7_valid_b(array_12_io_d_in_7_valid_b),
    .io_d_in_8_a(array_12_io_d_in_8_a),
    .io_d_in_8_valid_a(array_12_io_d_in_8_valid_a),
    .io_d_in_8_b(array_12_io_d_in_8_b),
    .io_d_in_8_valid_b(array_12_io_d_in_8_valid_b),
    .io_d_in_9_a(array_12_io_d_in_9_a),
    .io_d_in_9_valid_a(array_12_io_d_in_9_valid_a),
    .io_d_in_9_b(array_12_io_d_in_9_b),
    .io_d_in_9_valid_b(array_12_io_d_in_9_valid_b),
    .io_d_in_10_a(array_12_io_d_in_10_a),
    .io_d_in_10_valid_a(array_12_io_d_in_10_valid_a),
    .io_d_in_10_b(array_12_io_d_in_10_b),
    .io_d_in_10_valid_b(array_12_io_d_in_10_valid_b),
    .io_d_in_11_a(array_12_io_d_in_11_a),
    .io_d_in_11_valid_a(array_12_io_d_in_11_valid_a),
    .io_d_in_11_b(array_12_io_d_in_11_b),
    .io_d_in_11_valid_b(array_12_io_d_in_11_valid_b),
    .io_d_in_12_a(array_12_io_d_in_12_a),
    .io_d_in_12_valid_a(array_12_io_d_in_12_valid_a),
    .io_d_in_12_b(array_12_io_d_in_12_b),
    .io_d_in_12_valid_b(array_12_io_d_in_12_valid_b),
    .io_d_in_13_a(array_12_io_d_in_13_a),
    .io_d_in_13_valid_a(array_12_io_d_in_13_valid_a),
    .io_d_in_13_b(array_12_io_d_in_13_b),
    .io_d_in_13_valid_b(array_12_io_d_in_13_valid_b),
    .io_d_in_14_a(array_12_io_d_in_14_a),
    .io_d_in_14_valid_a(array_12_io_d_in_14_valid_a),
    .io_d_in_14_b(array_12_io_d_in_14_b),
    .io_d_in_14_valid_b(array_12_io_d_in_14_valid_b),
    .io_d_in_15_a(array_12_io_d_in_15_a),
    .io_d_in_15_valid_a(array_12_io_d_in_15_valid_a),
    .io_d_in_15_b(array_12_io_d_in_15_b),
    .io_d_in_15_valid_b(array_12_io_d_in_15_valid_b),
    .io_d_in_16_a(array_12_io_d_in_16_a),
    .io_d_in_16_valid_a(array_12_io_d_in_16_valid_a),
    .io_d_in_16_b(array_12_io_d_in_16_b),
    .io_d_in_16_valid_b(array_12_io_d_in_16_valid_b),
    .io_d_in_17_a(array_12_io_d_in_17_a),
    .io_d_in_17_valid_a(array_12_io_d_in_17_valid_a),
    .io_d_in_17_b(array_12_io_d_in_17_b),
    .io_d_in_17_valid_b(array_12_io_d_in_17_valid_b),
    .io_d_in_18_a(array_12_io_d_in_18_a),
    .io_d_in_18_valid_a(array_12_io_d_in_18_valid_a),
    .io_d_in_18_b(array_12_io_d_in_18_b),
    .io_d_in_18_valid_b(array_12_io_d_in_18_valid_b),
    .io_d_in_19_a(array_12_io_d_in_19_a),
    .io_d_in_19_valid_a(array_12_io_d_in_19_valid_a),
    .io_d_in_19_b(array_12_io_d_in_19_b),
    .io_d_in_19_valid_b(array_12_io_d_in_19_valid_b),
    .io_d_in_20_a(array_12_io_d_in_20_a),
    .io_d_in_20_valid_a(array_12_io_d_in_20_valid_a),
    .io_d_in_20_b(array_12_io_d_in_20_b),
    .io_d_in_20_valid_b(array_12_io_d_in_20_valid_b),
    .io_d_in_21_a(array_12_io_d_in_21_a),
    .io_d_in_21_valid_a(array_12_io_d_in_21_valid_a),
    .io_d_in_21_b(array_12_io_d_in_21_b),
    .io_d_in_21_valid_b(array_12_io_d_in_21_valid_b),
    .io_d_in_22_a(array_12_io_d_in_22_a),
    .io_d_in_22_valid_a(array_12_io_d_in_22_valid_a),
    .io_d_in_22_b(array_12_io_d_in_22_b),
    .io_d_in_22_valid_b(array_12_io_d_in_22_valid_b),
    .io_d_in_23_a(array_12_io_d_in_23_a),
    .io_d_in_23_valid_a(array_12_io_d_in_23_valid_a),
    .io_d_in_23_b(array_12_io_d_in_23_b),
    .io_d_in_23_valid_b(array_12_io_d_in_23_valid_b),
    .io_d_in_24_a(array_12_io_d_in_24_a),
    .io_d_in_24_valid_a(array_12_io_d_in_24_valid_a),
    .io_d_in_24_b(array_12_io_d_in_24_b),
    .io_d_in_24_valid_b(array_12_io_d_in_24_valid_b),
    .io_d_in_25_a(array_12_io_d_in_25_a),
    .io_d_in_25_valid_a(array_12_io_d_in_25_valid_a),
    .io_d_in_25_b(array_12_io_d_in_25_b),
    .io_d_in_25_valid_b(array_12_io_d_in_25_valid_b),
    .io_d_in_26_a(array_12_io_d_in_26_a),
    .io_d_in_26_valid_a(array_12_io_d_in_26_valid_a),
    .io_d_in_26_b(array_12_io_d_in_26_b),
    .io_d_in_26_valid_b(array_12_io_d_in_26_valid_b),
    .io_d_in_27_a(array_12_io_d_in_27_a),
    .io_d_in_27_valid_a(array_12_io_d_in_27_valid_a),
    .io_d_in_27_b(array_12_io_d_in_27_b),
    .io_d_in_27_valid_b(array_12_io_d_in_27_valid_b),
    .io_d_in_28_a(array_12_io_d_in_28_a),
    .io_d_in_28_valid_a(array_12_io_d_in_28_valid_a),
    .io_d_in_28_b(array_12_io_d_in_28_b),
    .io_d_in_28_valid_b(array_12_io_d_in_28_valid_b),
    .io_d_in_29_a(array_12_io_d_in_29_a),
    .io_d_in_29_valid_a(array_12_io_d_in_29_valid_a),
    .io_d_in_29_b(array_12_io_d_in_29_b),
    .io_d_in_29_valid_b(array_12_io_d_in_29_valid_b),
    .io_d_in_30_a(array_12_io_d_in_30_a),
    .io_d_in_30_valid_a(array_12_io_d_in_30_valid_a),
    .io_d_in_30_b(array_12_io_d_in_30_b),
    .io_d_in_30_valid_b(array_12_io_d_in_30_valid_b),
    .io_d_in_31_a(array_12_io_d_in_31_a),
    .io_d_in_31_valid_a(array_12_io_d_in_31_valid_a),
    .io_d_in_31_b(array_12_io_d_in_31_b),
    .io_d_in_31_valid_b(array_12_io_d_in_31_valid_b),
    .io_d_out_0_a(array_12_io_d_out_0_a),
    .io_d_out_0_valid_a(array_12_io_d_out_0_valid_a),
    .io_d_out_0_b(array_12_io_d_out_0_b),
    .io_d_out_0_valid_b(array_12_io_d_out_0_valid_b),
    .io_d_out_1_a(array_12_io_d_out_1_a),
    .io_d_out_1_valid_a(array_12_io_d_out_1_valid_a),
    .io_d_out_1_b(array_12_io_d_out_1_b),
    .io_d_out_1_valid_b(array_12_io_d_out_1_valid_b),
    .io_d_out_2_a(array_12_io_d_out_2_a),
    .io_d_out_2_valid_a(array_12_io_d_out_2_valid_a),
    .io_d_out_2_b(array_12_io_d_out_2_b),
    .io_d_out_2_valid_b(array_12_io_d_out_2_valid_b),
    .io_d_out_3_a(array_12_io_d_out_3_a),
    .io_d_out_3_valid_a(array_12_io_d_out_3_valid_a),
    .io_d_out_3_b(array_12_io_d_out_3_b),
    .io_d_out_3_valid_b(array_12_io_d_out_3_valid_b),
    .io_d_out_4_a(array_12_io_d_out_4_a),
    .io_d_out_4_valid_a(array_12_io_d_out_4_valid_a),
    .io_d_out_4_b(array_12_io_d_out_4_b),
    .io_d_out_4_valid_b(array_12_io_d_out_4_valid_b),
    .io_d_out_5_a(array_12_io_d_out_5_a),
    .io_d_out_5_valid_a(array_12_io_d_out_5_valid_a),
    .io_d_out_5_b(array_12_io_d_out_5_b),
    .io_d_out_5_valid_b(array_12_io_d_out_5_valid_b),
    .io_d_out_6_a(array_12_io_d_out_6_a),
    .io_d_out_6_valid_a(array_12_io_d_out_6_valid_a),
    .io_d_out_6_b(array_12_io_d_out_6_b),
    .io_d_out_6_valid_b(array_12_io_d_out_6_valid_b),
    .io_d_out_7_a(array_12_io_d_out_7_a),
    .io_d_out_7_valid_a(array_12_io_d_out_7_valid_a),
    .io_d_out_7_b(array_12_io_d_out_7_b),
    .io_d_out_7_valid_b(array_12_io_d_out_7_valid_b),
    .io_d_out_8_a(array_12_io_d_out_8_a),
    .io_d_out_8_valid_a(array_12_io_d_out_8_valid_a),
    .io_d_out_8_b(array_12_io_d_out_8_b),
    .io_d_out_8_valid_b(array_12_io_d_out_8_valid_b),
    .io_d_out_9_a(array_12_io_d_out_9_a),
    .io_d_out_9_valid_a(array_12_io_d_out_9_valid_a),
    .io_d_out_9_b(array_12_io_d_out_9_b),
    .io_d_out_9_valid_b(array_12_io_d_out_9_valid_b),
    .io_d_out_10_a(array_12_io_d_out_10_a),
    .io_d_out_10_valid_a(array_12_io_d_out_10_valid_a),
    .io_d_out_10_b(array_12_io_d_out_10_b),
    .io_d_out_10_valid_b(array_12_io_d_out_10_valid_b),
    .io_d_out_11_a(array_12_io_d_out_11_a),
    .io_d_out_11_valid_a(array_12_io_d_out_11_valid_a),
    .io_d_out_11_b(array_12_io_d_out_11_b),
    .io_d_out_11_valid_b(array_12_io_d_out_11_valid_b),
    .io_d_out_12_a(array_12_io_d_out_12_a),
    .io_d_out_12_valid_a(array_12_io_d_out_12_valid_a),
    .io_d_out_12_b(array_12_io_d_out_12_b),
    .io_d_out_12_valid_b(array_12_io_d_out_12_valid_b),
    .io_d_out_13_a(array_12_io_d_out_13_a),
    .io_d_out_13_valid_a(array_12_io_d_out_13_valid_a),
    .io_d_out_13_b(array_12_io_d_out_13_b),
    .io_d_out_13_valid_b(array_12_io_d_out_13_valid_b),
    .io_d_out_14_a(array_12_io_d_out_14_a),
    .io_d_out_14_valid_a(array_12_io_d_out_14_valid_a),
    .io_d_out_14_b(array_12_io_d_out_14_b),
    .io_d_out_14_valid_b(array_12_io_d_out_14_valid_b),
    .io_d_out_15_a(array_12_io_d_out_15_a),
    .io_d_out_15_valid_a(array_12_io_d_out_15_valid_a),
    .io_d_out_15_b(array_12_io_d_out_15_b),
    .io_d_out_15_valid_b(array_12_io_d_out_15_valid_b),
    .io_d_out_16_a(array_12_io_d_out_16_a),
    .io_d_out_16_valid_a(array_12_io_d_out_16_valid_a),
    .io_d_out_16_b(array_12_io_d_out_16_b),
    .io_d_out_16_valid_b(array_12_io_d_out_16_valid_b),
    .io_d_out_17_a(array_12_io_d_out_17_a),
    .io_d_out_17_valid_a(array_12_io_d_out_17_valid_a),
    .io_d_out_17_b(array_12_io_d_out_17_b),
    .io_d_out_17_valid_b(array_12_io_d_out_17_valid_b),
    .io_d_out_18_a(array_12_io_d_out_18_a),
    .io_d_out_18_valid_a(array_12_io_d_out_18_valid_a),
    .io_d_out_18_b(array_12_io_d_out_18_b),
    .io_d_out_18_valid_b(array_12_io_d_out_18_valid_b),
    .io_d_out_19_a(array_12_io_d_out_19_a),
    .io_d_out_19_valid_a(array_12_io_d_out_19_valid_a),
    .io_d_out_19_b(array_12_io_d_out_19_b),
    .io_d_out_19_valid_b(array_12_io_d_out_19_valid_b),
    .io_d_out_20_a(array_12_io_d_out_20_a),
    .io_d_out_20_valid_a(array_12_io_d_out_20_valid_a),
    .io_d_out_20_b(array_12_io_d_out_20_b),
    .io_d_out_20_valid_b(array_12_io_d_out_20_valid_b),
    .io_d_out_21_a(array_12_io_d_out_21_a),
    .io_d_out_21_valid_a(array_12_io_d_out_21_valid_a),
    .io_d_out_21_b(array_12_io_d_out_21_b),
    .io_d_out_21_valid_b(array_12_io_d_out_21_valid_b),
    .io_d_out_22_a(array_12_io_d_out_22_a),
    .io_d_out_22_valid_a(array_12_io_d_out_22_valid_a),
    .io_d_out_22_b(array_12_io_d_out_22_b),
    .io_d_out_22_valid_b(array_12_io_d_out_22_valid_b),
    .io_d_out_23_a(array_12_io_d_out_23_a),
    .io_d_out_23_valid_a(array_12_io_d_out_23_valid_a),
    .io_d_out_23_b(array_12_io_d_out_23_b),
    .io_d_out_23_valid_b(array_12_io_d_out_23_valid_b),
    .io_d_out_24_a(array_12_io_d_out_24_a),
    .io_d_out_24_valid_a(array_12_io_d_out_24_valid_a),
    .io_d_out_24_b(array_12_io_d_out_24_b),
    .io_d_out_24_valid_b(array_12_io_d_out_24_valid_b),
    .io_d_out_25_a(array_12_io_d_out_25_a),
    .io_d_out_25_valid_a(array_12_io_d_out_25_valid_a),
    .io_d_out_25_b(array_12_io_d_out_25_b),
    .io_d_out_25_valid_b(array_12_io_d_out_25_valid_b),
    .io_d_out_26_a(array_12_io_d_out_26_a),
    .io_d_out_26_valid_a(array_12_io_d_out_26_valid_a),
    .io_d_out_26_b(array_12_io_d_out_26_b),
    .io_d_out_26_valid_b(array_12_io_d_out_26_valid_b),
    .io_d_out_27_a(array_12_io_d_out_27_a),
    .io_d_out_27_valid_a(array_12_io_d_out_27_valid_a),
    .io_d_out_27_b(array_12_io_d_out_27_b),
    .io_d_out_27_valid_b(array_12_io_d_out_27_valid_b),
    .io_d_out_28_a(array_12_io_d_out_28_a),
    .io_d_out_28_valid_a(array_12_io_d_out_28_valid_a),
    .io_d_out_28_b(array_12_io_d_out_28_b),
    .io_d_out_28_valid_b(array_12_io_d_out_28_valid_b),
    .io_d_out_29_a(array_12_io_d_out_29_a),
    .io_d_out_29_valid_a(array_12_io_d_out_29_valid_a),
    .io_d_out_29_b(array_12_io_d_out_29_b),
    .io_d_out_29_valid_b(array_12_io_d_out_29_valid_b),
    .io_d_out_30_a(array_12_io_d_out_30_a),
    .io_d_out_30_valid_a(array_12_io_d_out_30_valid_a),
    .io_d_out_30_b(array_12_io_d_out_30_b),
    .io_d_out_30_valid_b(array_12_io_d_out_30_valid_b),
    .io_d_out_31_a(array_12_io_d_out_31_a),
    .io_d_out_31_valid_a(array_12_io_d_out_31_valid_a),
    .io_d_out_31_b(array_12_io_d_out_31_b),
    .io_d_out_31_valid_b(array_12_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_12_io_wr_en_mem1),
    .io_wr_en_mem2(array_12_io_wr_en_mem2),
    .io_wr_en_mem3(array_12_io_wr_en_mem3),
    .io_wr_en_mem4(array_12_io_wr_en_mem4),
    .io_wr_en_mem5(array_12_io_wr_en_mem5),
    .io_wr_en_mem6(array_12_io_wr_en_mem6),
    .io_wr_instr_mem1(array_12_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_12_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_12_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_12_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_12_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_12_io_wr_instr_mem6),
    .io_PC1_in(array_12_io_PC1_in),
    .io_PC6_out(array_12_io_PC6_out),
    .io_Addr_in(array_12_io_Addr_in),
    .io_Addr_out(array_12_io_Addr_out)
  );
  BuildingBlockNew array_13 ( // @[BP.scala 45:51]
    .clock(array_13_clock),
    .reset(array_13_reset),
    .io_d_in_0_a(array_13_io_d_in_0_a),
    .io_d_in_0_valid_a(array_13_io_d_in_0_valid_a),
    .io_d_in_0_b(array_13_io_d_in_0_b),
    .io_d_in_0_valid_b(array_13_io_d_in_0_valid_b),
    .io_d_in_1_a(array_13_io_d_in_1_a),
    .io_d_in_1_valid_a(array_13_io_d_in_1_valid_a),
    .io_d_in_1_b(array_13_io_d_in_1_b),
    .io_d_in_1_valid_b(array_13_io_d_in_1_valid_b),
    .io_d_in_2_a(array_13_io_d_in_2_a),
    .io_d_in_2_valid_a(array_13_io_d_in_2_valid_a),
    .io_d_in_2_b(array_13_io_d_in_2_b),
    .io_d_in_2_valid_b(array_13_io_d_in_2_valid_b),
    .io_d_in_3_a(array_13_io_d_in_3_a),
    .io_d_in_3_valid_a(array_13_io_d_in_3_valid_a),
    .io_d_in_3_b(array_13_io_d_in_3_b),
    .io_d_in_3_valid_b(array_13_io_d_in_3_valid_b),
    .io_d_in_4_a(array_13_io_d_in_4_a),
    .io_d_in_4_valid_a(array_13_io_d_in_4_valid_a),
    .io_d_in_4_b(array_13_io_d_in_4_b),
    .io_d_in_4_valid_b(array_13_io_d_in_4_valid_b),
    .io_d_in_5_a(array_13_io_d_in_5_a),
    .io_d_in_5_valid_a(array_13_io_d_in_5_valid_a),
    .io_d_in_5_b(array_13_io_d_in_5_b),
    .io_d_in_5_valid_b(array_13_io_d_in_5_valid_b),
    .io_d_in_6_a(array_13_io_d_in_6_a),
    .io_d_in_6_valid_a(array_13_io_d_in_6_valid_a),
    .io_d_in_6_b(array_13_io_d_in_6_b),
    .io_d_in_6_valid_b(array_13_io_d_in_6_valid_b),
    .io_d_in_7_a(array_13_io_d_in_7_a),
    .io_d_in_7_valid_a(array_13_io_d_in_7_valid_a),
    .io_d_in_7_b(array_13_io_d_in_7_b),
    .io_d_in_7_valid_b(array_13_io_d_in_7_valid_b),
    .io_d_in_8_a(array_13_io_d_in_8_a),
    .io_d_in_8_valid_a(array_13_io_d_in_8_valid_a),
    .io_d_in_8_b(array_13_io_d_in_8_b),
    .io_d_in_8_valid_b(array_13_io_d_in_8_valid_b),
    .io_d_in_9_a(array_13_io_d_in_9_a),
    .io_d_in_9_valid_a(array_13_io_d_in_9_valid_a),
    .io_d_in_9_b(array_13_io_d_in_9_b),
    .io_d_in_9_valid_b(array_13_io_d_in_9_valid_b),
    .io_d_in_10_a(array_13_io_d_in_10_a),
    .io_d_in_10_valid_a(array_13_io_d_in_10_valid_a),
    .io_d_in_10_b(array_13_io_d_in_10_b),
    .io_d_in_10_valid_b(array_13_io_d_in_10_valid_b),
    .io_d_in_11_a(array_13_io_d_in_11_a),
    .io_d_in_11_valid_a(array_13_io_d_in_11_valid_a),
    .io_d_in_11_b(array_13_io_d_in_11_b),
    .io_d_in_11_valid_b(array_13_io_d_in_11_valid_b),
    .io_d_in_12_a(array_13_io_d_in_12_a),
    .io_d_in_12_valid_a(array_13_io_d_in_12_valid_a),
    .io_d_in_12_b(array_13_io_d_in_12_b),
    .io_d_in_12_valid_b(array_13_io_d_in_12_valid_b),
    .io_d_in_13_a(array_13_io_d_in_13_a),
    .io_d_in_13_valid_a(array_13_io_d_in_13_valid_a),
    .io_d_in_13_b(array_13_io_d_in_13_b),
    .io_d_in_13_valid_b(array_13_io_d_in_13_valid_b),
    .io_d_in_14_a(array_13_io_d_in_14_a),
    .io_d_in_14_valid_a(array_13_io_d_in_14_valid_a),
    .io_d_in_14_b(array_13_io_d_in_14_b),
    .io_d_in_14_valid_b(array_13_io_d_in_14_valid_b),
    .io_d_in_15_a(array_13_io_d_in_15_a),
    .io_d_in_15_valid_a(array_13_io_d_in_15_valid_a),
    .io_d_in_15_b(array_13_io_d_in_15_b),
    .io_d_in_15_valid_b(array_13_io_d_in_15_valid_b),
    .io_d_in_16_a(array_13_io_d_in_16_a),
    .io_d_in_16_valid_a(array_13_io_d_in_16_valid_a),
    .io_d_in_16_b(array_13_io_d_in_16_b),
    .io_d_in_16_valid_b(array_13_io_d_in_16_valid_b),
    .io_d_in_17_a(array_13_io_d_in_17_a),
    .io_d_in_17_valid_a(array_13_io_d_in_17_valid_a),
    .io_d_in_17_b(array_13_io_d_in_17_b),
    .io_d_in_17_valid_b(array_13_io_d_in_17_valid_b),
    .io_d_in_18_a(array_13_io_d_in_18_a),
    .io_d_in_18_valid_a(array_13_io_d_in_18_valid_a),
    .io_d_in_18_b(array_13_io_d_in_18_b),
    .io_d_in_18_valid_b(array_13_io_d_in_18_valid_b),
    .io_d_in_19_a(array_13_io_d_in_19_a),
    .io_d_in_19_valid_a(array_13_io_d_in_19_valid_a),
    .io_d_in_19_b(array_13_io_d_in_19_b),
    .io_d_in_19_valid_b(array_13_io_d_in_19_valid_b),
    .io_d_in_20_a(array_13_io_d_in_20_a),
    .io_d_in_20_valid_a(array_13_io_d_in_20_valid_a),
    .io_d_in_20_b(array_13_io_d_in_20_b),
    .io_d_in_20_valid_b(array_13_io_d_in_20_valid_b),
    .io_d_in_21_a(array_13_io_d_in_21_a),
    .io_d_in_21_valid_a(array_13_io_d_in_21_valid_a),
    .io_d_in_21_b(array_13_io_d_in_21_b),
    .io_d_in_21_valid_b(array_13_io_d_in_21_valid_b),
    .io_d_in_22_a(array_13_io_d_in_22_a),
    .io_d_in_22_valid_a(array_13_io_d_in_22_valid_a),
    .io_d_in_22_b(array_13_io_d_in_22_b),
    .io_d_in_22_valid_b(array_13_io_d_in_22_valid_b),
    .io_d_in_23_a(array_13_io_d_in_23_a),
    .io_d_in_23_valid_a(array_13_io_d_in_23_valid_a),
    .io_d_in_23_b(array_13_io_d_in_23_b),
    .io_d_in_23_valid_b(array_13_io_d_in_23_valid_b),
    .io_d_in_24_a(array_13_io_d_in_24_a),
    .io_d_in_24_valid_a(array_13_io_d_in_24_valid_a),
    .io_d_in_24_b(array_13_io_d_in_24_b),
    .io_d_in_24_valid_b(array_13_io_d_in_24_valid_b),
    .io_d_in_25_a(array_13_io_d_in_25_a),
    .io_d_in_25_valid_a(array_13_io_d_in_25_valid_a),
    .io_d_in_25_b(array_13_io_d_in_25_b),
    .io_d_in_25_valid_b(array_13_io_d_in_25_valid_b),
    .io_d_in_26_a(array_13_io_d_in_26_a),
    .io_d_in_26_valid_a(array_13_io_d_in_26_valid_a),
    .io_d_in_26_b(array_13_io_d_in_26_b),
    .io_d_in_26_valid_b(array_13_io_d_in_26_valid_b),
    .io_d_in_27_a(array_13_io_d_in_27_a),
    .io_d_in_27_valid_a(array_13_io_d_in_27_valid_a),
    .io_d_in_27_b(array_13_io_d_in_27_b),
    .io_d_in_27_valid_b(array_13_io_d_in_27_valid_b),
    .io_d_in_28_a(array_13_io_d_in_28_a),
    .io_d_in_28_valid_a(array_13_io_d_in_28_valid_a),
    .io_d_in_28_b(array_13_io_d_in_28_b),
    .io_d_in_28_valid_b(array_13_io_d_in_28_valid_b),
    .io_d_in_29_a(array_13_io_d_in_29_a),
    .io_d_in_29_valid_a(array_13_io_d_in_29_valid_a),
    .io_d_in_29_b(array_13_io_d_in_29_b),
    .io_d_in_29_valid_b(array_13_io_d_in_29_valid_b),
    .io_d_in_30_a(array_13_io_d_in_30_a),
    .io_d_in_30_valid_a(array_13_io_d_in_30_valid_a),
    .io_d_in_30_b(array_13_io_d_in_30_b),
    .io_d_in_30_valid_b(array_13_io_d_in_30_valid_b),
    .io_d_in_31_a(array_13_io_d_in_31_a),
    .io_d_in_31_valid_a(array_13_io_d_in_31_valid_a),
    .io_d_in_31_b(array_13_io_d_in_31_b),
    .io_d_in_31_valid_b(array_13_io_d_in_31_valid_b),
    .io_d_out_0_a(array_13_io_d_out_0_a),
    .io_d_out_0_valid_a(array_13_io_d_out_0_valid_a),
    .io_d_out_0_b(array_13_io_d_out_0_b),
    .io_d_out_0_valid_b(array_13_io_d_out_0_valid_b),
    .io_d_out_1_a(array_13_io_d_out_1_a),
    .io_d_out_1_valid_a(array_13_io_d_out_1_valid_a),
    .io_d_out_1_b(array_13_io_d_out_1_b),
    .io_d_out_1_valid_b(array_13_io_d_out_1_valid_b),
    .io_d_out_2_a(array_13_io_d_out_2_a),
    .io_d_out_2_valid_a(array_13_io_d_out_2_valid_a),
    .io_d_out_2_b(array_13_io_d_out_2_b),
    .io_d_out_2_valid_b(array_13_io_d_out_2_valid_b),
    .io_d_out_3_a(array_13_io_d_out_3_a),
    .io_d_out_3_valid_a(array_13_io_d_out_3_valid_a),
    .io_d_out_3_b(array_13_io_d_out_3_b),
    .io_d_out_3_valid_b(array_13_io_d_out_3_valid_b),
    .io_d_out_4_a(array_13_io_d_out_4_a),
    .io_d_out_4_valid_a(array_13_io_d_out_4_valid_a),
    .io_d_out_4_b(array_13_io_d_out_4_b),
    .io_d_out_4_valid_b(array_13_io_d_out_4_valid_b),
    .io_d_out_5_a(array_13_io_d_out_5_a),
    .io_d_out_5_valid_a(array_13_io_d_out_5_valid_a),
    .io_d_out_5_b(array_13_io_d_out_5_b),
    .io_d_out_5_valid_b(array_13_io_d_out_5_valid_b),
    .io_d_out_6_a(array_13_io_d_out_6_a),
    .io_d_out_6_valid_a(array_13_io_d_out_6_valid_a),
    .io_d_out_6_b(array_13_io_d_out_6_b),
    .io_d_out_6_valid_b(array_13_io_d_out_6_valid_b),
    .io_d_out_7_a(array_13_io_d_out_7_a),
    .io_d_out_7_valid_a(array_13_io_d_out_7_valid_a),
    .io_d_out_7_b(array_13_io_d_out_7_b),
    .io_d_out_7_valid_b(array_13_io_d_out_7_valid_b),
    .io_d_out_8_a(array_13_io_d_out_8_a),
    .io_d_out_8_valid_a(array_13_io_d_out_8_valid_a),
    .io_d_out_8_b(array_13_io_d_out_8_b),
    .io_d_out_8_valid_b(array_13_io_d_out_8_valid_b),
    .io_d_out_9_a(array_13_io_d_out_9_a),
    .io_d_out_9_valid_a(array_13_io_d_out_9_valid_a),
    .io_d_out_9_b(array_13_io_d_out_9_b),
    .io_d_out_9_valid_b(array_13_io_d_out_9_valid_b),
    .io_d_out_10_a(array_13_io_d_out_10_a),
    .io_d_out_10_valid_a(array_13_io_d_out_10_valid_a),
    .io_d_out_10_b(array_13_io_d_out_10_b),
    .io_d_out_10_valid_b(array_13_io_d_out_10_valid_b),
    .io_d_out_11_a(array_13_io_d_out_11_a),
    .io_d_out_11_valid_a(array_13_io_d_out_11_valid_a),
    .io_d_out_11_b(array_13_io_d_out_11_b),
    .io_d_out_11_valid_b(array_13_io_d_out_11_valid_b),
    .io_d_out_12_a(array_13_io_d_out_12_a),
    .io_d_out_12_valid_a(array_13_io_d_out_12_valid_a),
    .io_d_out_12_b(array_13_io_d_out_12_b),
    .io_d_out_12_valid_b(array_13_io_d_out_12_valid_b),
    .io_d_out_13_a(array_13_io_d_out_13_a),
    .io_d_out_13_valid_a(array_13_io_d_out_13_valid_a),
    .io_d_out_13_b(array_13_io_d_out_13_b),
    .io_d_out_13_valid_b(array_13_io_d_out_13_valid_b),
    .io_d_out_14_a(array_13_io_d_out_14_a),
    .io_d_out_14_valid_a(array_13_io_d_out_14_valid_a),
    .io_d_out_14_b(array_13_io_d_out_14_b),
    .io_d_out_14_valid_b(array_13_io_d_out_14_valid_b),
    .io_d_out_15_a(array_13_io_d_out_15_a),
    .io_d_out_15_valid_a(array_13_io_d_out_15_valid_a),
    .io_d_out_15_b(array_13_io_d_out_15_b),
    .io_d_out_15_valid_b(array_13_io_d_out_15_valid_b),
    .io_d_out_16_a(array_13_io_d_out_16_a),
    .io_d_out_16_valid_a(array_13_io_d_out_16_valid_a),
    .io_d_out_16_b(array_13_io_d_out_16_b),
    .io_d_out_16_valid_b(array_13_io_d_out_16_valid_b),
    .io_d_out_17_a(array_13_io_d_out_17_a),
    .io_d_out_17_valid_a(array_13_io_d_out_17_valid_a),
    .io_d_out_17_b(array_13_io_d_out_17_b),
    .io_d_out_17_valid_b(array_13_io_d_out_17_valid_b),
    .io_d_out_18_a(array_13_io_d_out_18_a),
    .io_d_out_18_valid_a(array_13_io_d_out_18_valid_a),
    .io_d_out_18_b(array_13_io_d_out_18_b),
    .io_d_out_18_valid_b(array_13_io_d_out_18_valid_b),
    .io_d_out_19_a(array_13_io_d_out_19_a),
    .io_d_out_19_valid_a(array_13_io_d_out_19_valid_a),
    .io_d_out_19_b(array_13_io_d_out_19_b),
    .io_d_out_19_valid_b(array_13_io_d_out_19_valid_b),
    .io_d_out_20_a(array_13_io_d_out_20_a),
    .io_d_out_20_valid_a(array_13_io_d_out_20_valid_a),
    .io_d_out_20_b(array_13_io_d_out_20_b),
    .io_d_out_20_valid_b(array_13_io_d_out_20_valid_b),
    .io_d_out_21_a(array_13_io_d_out_21_a),
    .io_d_out_21_valid_a(array_13_io_d_out_21_valid_a),
    .io_d_out_21_b(array_13_io_d_out_21_b),
    .io_d_out_21_valid_b(array_13_io_d_out_21_valid_b),
    .io_d_out_22_a(array_13_io_d_out_22_a),
    .io_d_out_22_valid_a(array_13_io_d_out_22_valid_a),
    .io_d_out_22_b(array_13_io_d_out_22_b),
    .io_d_out_22_valid_b(array_13_io_d_out_22_valid_b),
    .io_d_out_23_a(array_13_io_d_out_23_a),
    .io_d_out_23_valid_a(array_13_io_d_out_23_valid_a),
    .io_d_out_23_b(array_13_io_d_out_23_b),
    .io_d_out_23_valid_b(array_13_io_d_out_23_valid_b),
    .io_d_out_24_a(array_13_io_d_out_24_a),
    .io_d_out_24_valid_a(array_13_io_d_out_24_valid_a),
    .io_d_out_24_b(array_13_io_d_out_24_b),
    .io_d_out_24_valid_b(array_13_io_d_out_24_valid_b),
    .io_d_out_25_a(array_13_io_d_out_25_a),
    .io_d_out_25_valid_a(array_13_io_d_out_25_valid_a),
    .io_d_out_25_b(array_13_io_d_out_25_b),
    .io_d_out_25_valid_b(array_13_io_d_out_25_valid_b),
    .io_d_out_26_a(array_13_io_d_out_26_a),
    .io_d_out_26_valid_a(array_13_io_d_out_26_valid_a),
    .io_d_out_26_b(array_13_io_d_out_26_b),
    .io_d_out_26_valid_b(array_13_io_d_out_26_valid_b),
    .io_d_out_27_a(array_13_io_d_out_27_a),
    .io_d_out_27_valid_a(array_13_io_d_out_27_valid_a),
    .io_d_out_27_b(array_13_io_d_out_27_b),
    .io_d_out_27_valid_b(array_13_io_d_out_27_valid_b),
    .io_d_out_28_a(array_13_io_d_out_28_a),
    .io_d_out_28_valid_a(array_13_io_d_out_28_valid_a),
    .io_d_out_28_b(array_13_io_d_out_28_b),
    .io_d_out_28_valid_b(array_13_io_d_out_28_valid_b),
    .io_d_out_29_a(array_13_io_d_out_29_a),
    .io_d_out_29_valid_a(array_13_io_d_out_29_valid_a),
    .io_d_out_29_b(array_13_io_d_out_29_b),
    .io_d_out_29_valid_b(array_13_io_d_out_29_valid_b),
    .io_d_out_30_a(array_13_io_d_out_30_a),
    .io_d_out_30_valid_a(array_13_io_d_out_30_valid_a),
    .io_d_out_30_b(array_13_io_d_out_30_b),
    .io_d_out_30_valid_b(array_13_io_d_out_30_valid_b),
    .io_d_out_31_a(array_13_io_d_out_31_a),
    .io_d_out_31_valid_a(array_13_io_d_out_31_valid_a),
    .io_d_out_31_b(array_13_io_d_out_31_b),
    .io_d_out_31_valid_b(array_13_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_13_io_wr_en_mem1),
    .io_wr_en_mem2(array_13_io_wr_en_mem2),
    .io_wr_en_mem3(array_13_io_wr_en_mem3),
    .io_wr_en_mem4(array_13_io_wr_en_mem4),
    .io_wr_en_mem5(array_13_io_wr_en_mem5),
    .io_wr_en_mem6(array_13_io_wr_en_mem6),
    .io_wr_instr_mem1(array_13_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_13_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_13_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_13_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_13_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_13_io_wr_instr_mem6),
    .io_PC1_in(array_13_io_PC1_in),
    .io_PC6_out(array_13_io_PC6_out),
    .io_Addr_in(array_13_io_Addr_in),
    .io_Addr_out(array_13_io_Addr_out)
  );
  BuildingBlockNew array_14 ( // @[BP.scala 45:51]
    .clock(array_14_clock),
    .reset(array_14_reset),
    .io_d_in_0_a(array_14_io_d_in_0_a),
    .io_d_in_0_valid_a(array_14_io_d_in_0_valid_a),
    .io_d_in_0_b(array_14_io_d_in_0_b),
    .io_d_in_0_valid_b(array_14_io_d_in_0_valid_b),
    .io_d_in_1_a(array_14_io_d_in_1_a),
    .io_d_in_1_valid_a(array_14_io_d_in_1_valid_a),
    .io_d_in_1_b(array_14_io_d_in_1_b),
    .io_d_in_1_valid_b(array_14_io_d_in_1_valid_b),
    .io_d_in_2_a(array_14_io_d_in_2_a),
    .io_d_in_2_valid_a(array_14_io_d_in_2_valid_a),
    .io_d_in_2_b(array_14_io_d_in_2_b),
    .io_d_in_2_valid_b(array_14_io_d_in_2_valid_b),
    .io_d_in_3_a(array_14_io_d_in_3_a),
    .io_d_in_3_valid_a(array_14_io_d_in_3_valid_a),
    .io_d_in_3_b(array_14_io_d_in_3_b),
    .io_d_in_3_valid_b(array_14_io_d_in_3_valid_b),
    .io_d_in_4_a(array_14_io_d_in_4_a),
    .io_d_in_4_valid_a(array_14_io_d_in_4_valid_a),
    .io_d_in_4_b(array_14_io_d_in_4_b),
    .io_d_in_4_valid_b(array_14_io_d_in_4_valid_b),
    .io_d_in_5_a(array_14_io_d_in_5_a),
    .io_d_in_5_valid_a(array_14_io_d_in_5_valid_a),
    .io_d_in_5_b(array_14_io_d_in_5_b),
    .io_d_in_5_valid_b(array_14_io_d_in_5_valid_b),
    .io_d_in_6_a(array_14_io_d_in_6_a),
    .io_d_in_6_valid_a(array_14_io_d_in_6_valid_a),
    .io_d_in_6_b(array_14_io_d_in_6_b),
    .io_d_in_6_valid_b(array_14_io_d_in_6_valid_b),
    .io_d_in_7_a(array_14_io_d_in_7_a),
    .io_d_in_7_valid_a(array_14_io_d_in_7_valid_a),
    .io_d_in_7_b(array_14_io_d_in_7_b),
    .io_d_in_7_valid_b(array_14_io_d_in_7_valid_b),
    .io_d_in_8_a(array_14_io_d_in_8_a),
    .io_d_in_8_valid_a(array_14_io_d_in_8_valid_a),
    .io_d_in_8_b(array_14_io_d_in_8_b),
    .io_d_in_8_valid_b(array_14_io_d_in_8_valid_b),
    .io_d_in_9_a(array_14_io_d_in_9_a),
    .io_d_in_9_valid_a(array_14_io_d_in_9_valid_a),
    .io_d_in_9_b(array_14_io_d_in_9_b),
    .io_d_in_9_valid_b(array_14_io_d_in_9_valid_b),
    .io_d_in_10_a(array_14_io_d_in_10_a),
    .io_d_in_10_valid_a(array_14_io_d_in_10_valid_a),
    .io_d_in_10_b(array_14_io_d_in_10_b),
    .io_d_in_10_valid_b(array_14_io_d_in_10_valid_b),
    .io_d_in_11_a(array_14_io_d_in_11_a),
    .io_d_in_11_valid_a(array_14_io_d_in_11_valid_a),
    .io_d_in_11_b(array_14_io_d_in_11_b),
    .io_d_in_11_valid_b(array_14_io_d_in_11_valid_b),
    .io_d_in_12_a(array_14_io_d_in_12_a),
    .io_d_in_12_valid_a(array_14_io_d_in_12_valid_a),
    .io_d_in_12_b(array_14_io_d_in_12_b),
    .io_d_in_12_valid_b(array_14_io_d_in_12_valid_b),
    .io_d_in_13_a(array_14_io_d_in_13_a),
    .io_d_in_13_valid_a(array_14_io_d_in_13_valid_a),
    .io_d_in_13_b(array_14_io_d_in_13_b),
    .io_d_in_13_valid_b(array_14_io_d_in_13_valid_b),
    .io_d_in_14_a(array_14_io_d_in_14_a),
    .io_d_in_14_valid_a(array_14_io_d_in_14_valid_a),
    .io_d_in_14_b(array_14_io_d_in_14_b),
    .io_d_in_14_valid_b(array_14_io_d_in_14_valid_b),
    .io_d_in_15_a(array_14_io_d_in_15_a),
    .io_d_in_15_valid_a(array_14_io_d_in_15_valid_a),
    .io_d_in_15_b(array_14_io_d_in_15_b),
    .io_d_in_15_valid_b(array_14_io_d_in_15_valid_b),
    .io_d_in_16_a(array_14_io_d_in_16_a),
    .io_d_in_16_valid_a(array_14_io_d_in_16_valid_a),
    .io_d_in_16_b(array_14_io_d_in_16_b),
    .io_d_in_16_valid_b(array_14_io_d_in_16_valid_b),
    .io_d_in_17_a(array_14_io_d_in_17_a),
    .io_d_in_17_valid_a(array_14_io_d_in_17_valid_a),
    .io_d_in_17_b(array_14_io_d_in_17_b),
    .io_d_in_17_valid_b(array_14_io_d_in_17_valid_b),
    .io_d_in_18_a(array_14_io_d_in_18_a),
    .io_d_in_18_valid_a(array_14_io_d_in_18_valid_a),
    .io_d_in_18_b(array_14_io_d_in_18_b),
    .io_d_in_18_valid_b(array_14_io_d_in_18_valid_b),
    .io_d_in_19_a(array_14_io_d_in_19_a),
    .io_d_in_19_valid_a(array_14_io_d_in_19_valid_a),
    .io_d_in_19_b(array_14_io_d_in_19_b),
    .io_d_in_19_valid_b(array_14_io_d_in_19_valid_b),
    .io_d_in_20_a(array_14_io_d_in_20_a),
    .io_d_in_20_valid_a(array_14_io_d_in_20_valid_a),
    .io_d_in_20_b(array_14_io_d_in_20_b),
    .io_d_in_20_valid_b(array_14_io_d_in_20_valid_b),
    .io_d_in_21_a(array_14_io_d_in_21_a),
    .io_d_in_21_valid_a(array_14_io_d_in_21_valid_a),
    .io_d_in_21_b(array_14_io_d_in_21_b),
    .io_d_in_21_valid_b(array_14_io_d_in_21_valid_b),
    .io_d_in_22_a(array_14_io_d_in_22_a),
    .io_d_in_22_valid_a(array_14_io_d_in_22_valid_a),
    .io_d_in_22_b(array_14_io_d_in_22_b),
    .io_d_in_22_valid_b(array_14_io_d_in_22_valid_b),
    .io_d_in_23_a(array_14_io_d_in_23_a),
    .io_d_in_23_valid_a(array_14_io_d_in_23_valid_a),
    .io_d_in_23_b(array_14_io_d_in_23_b),
    .io_d_in_23_valid_b(array_14_io_d_in_23_valid_b),
    .io_d_in_24_a(array_14_io_d_in_24_a),
    .io_d_in_24_valid_a(array_14_io_d_in_24_valid_a),
    .io_d_in_24_b(array_14_io_d_in_24_b),
    .io_d_in_24_valid_b(array_14_io_d_in_24_valid_b),
    .io_d_in_25_a(array_14_io_d_in_25_a),
    .io_d_in_25_valid_a(array_14_io_d_in_25_valid_a),
    .io_d_in_25_b(array_14_io_d_in_25_b),
    .io_d_in_25_valid_b(array_14_io_d_in_25_valid_b),
    .io_d_in_26_a(array_14_io_d_in_26_a),
    .io_d_in_26_valid_a(array_14_io_d_in_26_valid_a),
    .io_d_in_26_b(array_14_io_d_in_26_b),
    .io_d_in_26_valid_b(array_14_io_d_in_26_valid_b),
    .io_d_in_27_a(array_14_io_d_in_27_a),
    .io_d_in_27_valid_a(array_14_io_d_in_27_valid_a),
    .io_d_in_27_b(array_14_io_d_in_27_b),
    .io_d_in_27_valid_b(array_14_io_d_in_27_valid_b),
    .io_d_in_28_a(array_14_io_d_in_28_a),
    .io_d_in_28_valid_a(array_14_io_d_in_28_valid_a),
    .io_d_in_28_b(array_14_io_d_in_28_b),
    .io_d_in_28_valid_b(array_14_io_d_in_28_valid_b),
    .io_d_in_29_a(array_14_io_d_in_29_a),
    .io_d_in_29_valid_a(array_14_io_d_in_29_valid_a),
    .io_d_in_29_b(array_14_io_d_in_29_b),
    .io_d_in_29_valid_b(array_14_io_d_in_29_valid_b),
    .io_d_in_30_a(array_14_io_d_in_30_a),
    .io_d_in_30_valid_a(array_14_io_d_in_30_valid_a),
    .io_d_in_30_b(array_14_io_d_in_30_b),
    .io_d_in_30_valid_b(array_14_io_d_in_30_valid_b),
    .io_d_in_31_a(array_14_io_d_in_31_a),
    .io_d_in_31_valid_a(array_14_io_d_in_31_valid_a),
    .io_d_in_31_b(array_14_io_d_in_31_b),
    .io_d_in_31_valid_b(array_14_io_d_in_31_valid_b),
    .io_d_out_0_a(array_14_io_d_out_0_a),
    .io_d_out_0_valid_a(array_14_io_d_out_0_valid_a),
    .io_d_out_0_b(array_14_io_d_out_0_b),
    .io_d_out_0_valid_b(array_14_io_d_out_0_valid_b),
    .io_d_out_1_a(array_14_io_d_out_1_a),
    .io_d_out_1_valid_a(array_14_io_d_out_1_valid_a),
    .io_d_out_1_b(array_14_io_d_out_1_b),
    .io_d_out_1_valid_b(array_14_io_d_out_1_valid_b),
    .io_d_out_2_a(array_14_io_d_out_2_a),
    .io_d_out_2_valid_a(array_14_io_d_out_2_valid_a),
    .io_d_out_2_b(array_14_io_d_out_2_b),
    .io_d_out_2_valid_b(array_14_io_d_out_2_valid_b),
    .io_d_out_3_a(array_14_io_d_out_3_a),
    .io_d_out_3_valid_a(array_14_io_d_out_3_valid_a),
    .io_d_out_3_b(array_14_io_d_out_3_b),
    .io_d_out_3_valid_b(array_14_io_d_out_3_valid_b),
    .io_d_out_4_a(array_14_io_d_out_4_a),
    .io_d_out_4_valid_a(array_14_io_d_out_4_valid_a),
    .io_d_out_4_b(array_14_io_d_out_4_b),
    .io_d_out_4_valid_b(array_14_io_d_out_4_valid_b),
    .io_d_out_5_a(array_14_io_d_out_5_a),
    .io_d_out_5_valid_a(array_14_io_d_out_5_valid_a),
    .io_d_out_5_b(array_14_io_d_out_5_b),
    .io_d_out_5_valid_b(array_14_io_d_out_5_valid_b),
    .io_d_out_6_a(array_14_io_d_out_6_a),
    .io_d_out_6_valid_a(array_14_io_d_out_6_valid_a),
    .io_d_out_6_b(array_14_io_d_out_6_b),
    .io_d_out_6_valid_b(array_14_io_d_out_6_valid_b),
    .io_d_out_7_a(array_14_io_d_out_7_a),
    .io_d_out_7_valid_a(array_14_io_d_out_7_valid_a),
    .io_d_out_7_b(array_14_io_d_out_7_b),
    .io_d_out_7_valid_b(array_14_io_d_out_7_valid_b),
    .io_d_out_8_a(array_14_io_d_out_8_a),
    .io_d_out_8_valid_a(array_14_io_d_out_8_valid_a),
    .io_d_out_8_b(array_14_io_d_out_8_b),
    .io_d_out_8_valid_b(array_14_io_d_out_8_valid_b),
    .io_d_out_9_a(array_14_io_d_out_9_a),
    .io_d_out_9_valid_a(array_14_io_d_out_9_valid_a),
    .io_d_out_9_b(array_14_io_d_out_9_b),
    .io_d_out_9_valid_b(array_14_io_d_out_9_valid_b),
    .io_d_out_10_a(array_14_io_d_out_10_a),
    .io_d_out_10_valid_a(array_14_io_d_out_10_valid_a),
    .io_d_out_10_b(array_14_io_d_out_10_b),
    .io_d_out_10_valid_b(array_14_io_d_out_10_valid_b),
    .io_d_out_11_a(array_14_io_d_out_11_a),
    .io_d_out_11_valid_a(array_14_io_d_out_11_valid_a),
    .io_d_out_11_b(array_14_io_d_out_11_b),
    .io_d_out_11_valid_b(array_14_io_d_out_11_valid_b),
    .io_d_out_12_a(array_14_io_d_out_12_a),
    .io_d_out_12_valid_a(array_14_io_d_out_12_valid_a),
    .io_d_out_12_b(array_14_io_d_out_12_b),
    .io_d_out_12_valid_b(array_14_io_d_out_12_valid_b),
    .io_d_out_13_a(array_14_io_d_out_13_a),
    .io_d_out_13_valid_a(array_14_io_d_out_13_valid_a),
    .io_d_out_13_b(array_14_io_d_out_13_b),
    .io_d_out_13_valid_b(array_14_io_d_out_13_valid_b),
    .io_d_out_14_a(array_14_io_d_out_14_a),
    .io_d_out_14_valid_a(array_14_io_d_out_14_valid_a),
    .io_d_out_14_b(array_14_io_d_out_14_b),
    .io_d_out_14_valid_b(array_14_io_d_out_14_valid_b),
    .io_d_out_15_a(array_14_io_d_out_15_a),
    .io_d_out_15_valid_a(array_14_io_d_out_15_valid_a),
    .io_d_out_15_b(array_14_io_d_out_15_b),
    .io_d_out_15_valid_b(array_14_io_d_out_15_valid_b),
    .io_d_out_16_a(array_14_io_d_out_16_a),
    .io_d_out_16_valid_a(array_14_io_d_out_16_valid_a),
    .io_d_out_16_b(array_14_io_d_out_16_b),
    .io_d_out_16_valid_b(array_14_io_d_out_16_valid_b),
    .io_d_out_17_a(array_14_io_d_out_17_a),
    .io_d_out_17_valid_a(array_14_io_d_out_17_valid_a),
    .io_d_out_17_b(array_14_io_d_out_17_b),
    .io_d_out_17_valid_b(array_14_io_d_out_17_valid_b),
    .io_d_out_18_a(array_14_io_d_out_18_a),
    .io_d_out_18_valid_a(array_14_io_d_out_18_valid_a),
    .io_d_out_18_b(array_14_io_d_out_18_b),
    .io_d_out_18_valid_b(array_14_io_d_out_18_valid_b),
    .io_d_out_19_a(array_14_io_d_out_19_a),
    .io_d_out_19_valid_a(array_14_io_d_out_19_valid_a),
    .io_d_out_19_b(array_14_io_d_out_19_b),
    .io_d_out_19_valid_b(array_14_io_d_out_19_valid_b),
    .io_d_out_20_a(array_14_io_d_out_20_a),
    .io_d_out_20_valid_a(array_14_io_d_out_20_valid_a),
    .io_d_out_20_b(array_14_io_d_out_20_b),
    .io_d_out_20_valid_b(array_14_io_d_out_20_valid_b),
    .io_d_out_21_a(array_14_io_d_out_21_a),
    .io_d_out_21_valid_a(array_14_io_d_out_21_valid_a),
    .io_d_out_21_b(array_14_io_d_out_21_b),
    .io_d_out_21_valid_b(array_14_io_d_out_21_valid_b),
    .io_d_out_22_a(array_14_io_d_out_22_a),
    .io_d_out_22_valid_a(array_14_io_d_out_22_valid_a),
    .io_d_out_22_b(array_14_io_d_out_22_b),
    .io_d_out_22_valid_b(array_14_io_d_out_22_valid_b),
    .io_d_out_23_a(array_14_io_d_out_23_a),
    .io_d_out_23_valid_a(array_14_io_d_out_23_valid_a),
    .io_d_out_23_b(array_14_io_d_out_23_b),
    .io_d_out_23_valid_b(array_14_io_d_out_23_valid_b),
    .io_d_out_24_a(array_14_io_d_out_24_a),
    .io_d_out_24_valid_a(array_14_io_d_out_24_valid_a),
    .io_d_out_24_b(array_14_io_d_out_24_b),
    .io_d_out_24_valid_b(array_14_io_d_out_24_valid_b),
    .io_d_out_25_a(array_14_io_d_out_25_a),
    .io_d_out_25_valid_a(array_14_io_d_out_25_valid_a),
    .io_d_out_25_b(array_14_io_d_out_25_b),
    .io_d_out_25_valid_b(array_14_io_d_out_25_valid_b),
    .io_d_out_26_a(array_14_io_d_out_26_a),
    .io_d_out_26_valid_a(array_14_io_d_out_26_valid_a),
    .io_d_out_26_b(array_14_io_d_out_26_b),
    .io_d_out_26_valid_b(array_14_io_d_out_26_valid_b),
    .io_d_out_27_a(array_14_io_d_out_27_a),
    .io_d_out_27_valid_a(array_14_io_d_out_27_valid_a),
    .io_d_out_27_b(array_14_io_d_out_27_b),
    .io_d_out_27_valid_b(array_14_io_d_out_27_valid_b),
    .io_d_out_28_a(array_14_io_d_out_28_a),
    .io_d_out_28_valid_a(array_14_io_d_out_28_valid_a),
    .io_d_out_28_b(array_14_io_d_out_28_b),
    .io_d_out_28_valid_b(array_14_io_d_out_28_valid_b),
    .io_d_out_29_a(array_14_io_d_out_29_a),
    .io_d_out_29_valid_a(array_14_io_d_out_29_valid_a),
    .io_d_out_29_b(array_14_io_d_out_29_b),
    .io_d_out_29_valid_b(array_14_io_d_out_29_valid_b),
    .io_d_out_30_a(array_14_io_d_out_30_a),
    .io_d_out_30_valid_a(array_14_io_d_out_30_valid_a),
    .io_d_out_30_b(array_14_io_d_out_30_b),
    .io_d_out_30_valid_b(array_14_io_d_out_30_valid_b),
    .io_d_out_31_a(array_14_io_d_out_31_a),
    .io_d_out_31_valid_a(array_14_io_d_out_31_valid_a),
    .io_d_out_31_b(array_14_io_d_out_31_b),
    .io_d_out_31_valid_b(array_14_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_14_io_wr_en_mem1),
    .io_wr_en_mem2(array_14_io_wr_en_mem2),
    .io_wr_en_mem3(array_14_io_wr_en_mem3),
    .io_wr_en_mem4(array_14_io_wr_en_mem4),
    .io_wr_en_mem5(array_14_io_wr_en_mem5),
    .io_wr_en_mem6(array_14_io_wr_en_mem6),
    .io_wr_instr_mem1(array_14_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_14_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_14_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_14_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_14_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_14_io_wr_instr_mem6),
    .io_PC1_in(array_14_io_PC1_in),
    .io_PC6_out(array_14_io_PC6_out),
    .io_Addr_in(array_14_io_Addr_in),
    .io_Addr_out(array_14_io_Addr_out)
  );
  BuildingBlockNew array_15 ( // @[BP.scala 45:51]
    .clock(array_15_clock),
    .reset(array_15_reset),
    .io_d_in_0_a(array_15_io_d_in_0_a),
    .io_d_in_0_valid_a(array_15_io_d_in_0_valid_a),
    .io_d_in_0_b(array_15_io_d_in_0_b),
    .io_d_in_0_valid_b(array_15_io_d_in_0_valid_b),
    .io_d_in_1_a(array_15_io_d_in_1_a),
    .io_d_in_1_valid_a(array_15_io_d_in_1_valid_a),
    .io_d_in_1_b(array_15_io_d_in_1_b),
    .io_d_in_1_valid_b(array_15_io_d_in_1_valid_b),
    .io_d_in_2_a(array_15_io_d_in_2_a),
    .io_d_in_2_valid_a(array_15_io_d_in_2_valid_a),
    .io_d_in_2_b(array_15_io_d_in_2_b),
    .io_d_in_2_valid_b(array_15_io_d_in_2_valid_b),
    .io_d_in_3_a(array_15_io_d_in_3_a),
    .io_d_in_3_valid_a(array_15_io_d_in_3_valid_a),
    .io_d_in_3_b(array_15_io_d_in_3_b),
    .io_d_in_3_valid_b(array_15_io_d_in_3_valid_b),
    .io_d_in_4_a(array_15_io_d_in_4_a),
    .io_d_in_4_valid_a(array_15_io_d_in_4_valid_a),
    .io_d_in_4_b(array_15_io_d_in_4_b),
    .io_d_in_4_valid_b(array_15_io_d_in_4_valid_b),
    .io_d_in_5_a(array_15_io_d_in_5_a),
    .io_d_in_5_valid_a(array_15_io_d_in_5_valid_a),
    .io_d_in_5_b(array_15_io_d_in_5_b),
    .io_d_in_5_valid_b(array_15_io_d_in_5_valid_b),
    .io_d_in_6_a(array_15_io_d_in_6_a),
    .io_d_in_6_valid_a(array_15_io_d_in_6_valid_a),
    .io_d_in_6_b(array_15_io_d_in_6_b),
    .io_d_in_6_valid_b(array_15_io_d_in_6_valid_b),
    .io_d_in_7_a(array_15_io_d_in_7_a),
    .io_d_in_7_valid_a(array_15_io_d_in_7_valid_a),
    .io_d_in_7_b(array_15_io_d_in_7_b),
    .io_d_in_7_valid_b(array_15_io_d_in_7_valid_b),
    .io_d_in_8_a(array_15_io_d_in_8_a),
    .io_d_in_8_valid_a(array_15_io_d_in_8_valid_a),
    .io_d_in_8_b(array_15_io_d_in_8_b),
    .io_d_in_8_valid_b(array_15_io_d_in_8_valid_b),
    .io_d_in_9_a(array_15_io_d_in_9_a),
    .io_d_in_9_valid_a(array_15_io_d_in_9_valid_a),
    .io_d_in_9_b(array_15_io_d_in_9_b),
    .io_d_in_9_valid_b(array_15_io_d_in_9_valid_b),
    .io_d_in_10_a(array_15_io_d_in_10_a),
    .io_d_in_10_valid_a(array_15_io_d_in_10_valid_a),
    .io_d_in_10_b(array_15_io_d_in_10_b),
    .io_d_in_10_valid_b(array_15_io_d_in_10_valid_b),
    .io_d_in_11_a(array_15_io_d_in_11_a),
    .io_d_in_11_valid_a(array_15_io_d_in_11_valid_a),
    .io_d_in_11_b(array_15_io_d_in_11_b),
    .io_d_in_11_valid_b(array_15_io_d_in_11_valid_b),
    .io_d_in_12_a(array_15_io_d_in_12_a),
    .io_d_in_12_valid_a(array_15_io_d_in_12_valid_a),
    .io_d_in_12_b(array_15_io_d_in_12_b),
    .io_d_in_12_valid_b(array_15_io_d_in_12_valid_b),
    .io_d_in_13_a(array_15_io_d_in_13_a),
    .io_d_in_13_valid_a(array_15_io_d_in_13_valid_a),
    .io_d_in_13_b(array_15_io_d_in_13_b),
    .io_d_in_13_valid_b(array_15_io_d_in_13_valid_b),
    .io_d_in_14_a(array_15_io_d_in_14_a),
    .io_d_in_14_valid_a(array_15_io_d_in_14_valid_a),
    .io_d_in_14_b(array_15_io_d_in_14_b),
    .io_d_in_14_valid_b(array_15_io_d_in_14_valid_b),
    .io_d_in_15_a(array_15_io_d_in_15_a),
    .io_d_in_15_valid_a(array_15_io_d_in_15_valid_a),
    .io_d_in_15_b(array_15_io_d_in_15_b),
    .io_d_in_15_valid_b(array_15_io_d_in_15_valid_b),
    .io_d_in_16_a(array_15_io_d_in_16_a),
    .io_d_in_16_valid_a(array_15_io_d_in_16_valid_a),
    .io_d_in_16_b(array_15_io_d_in_16_b),
    .io_d_in_16_valid_b(array_15_io_d_in_16_valid_b),
    .io_d_in_17_a(array_15_io_d_in_17_a),
    .io_d_in_17_valid_a(array_15_io_d_in_17_valid_a),
    .io_d_in_17_b(array_15_io_d_in_17_b),
    .io_d_in_17_valid_b(array_15_io_d_in_17_valid_b),
    .io_d_in_18_a(array_15_io_d_in_18_a),
    .io_d_in_18_valid_a(array_15_io_d_in_18_valid_a),
    .io_d_in_18_b(array_15_io_d_in_18_b),
    .io_d_in_18_valid_b(array_15_io_d_in_18_valid_b),
    .io_d_in_19_a(array_15_io_d_in_19_a),
    .io_d_in_19_valid_a(array_15_io_d_in_19_valid_a),
    .io_d_in_19_b(array_15_io_d_in_19_b),
    .io_d_in_19_valid_b(array_15_io_d_in_19_valid_b),
    .io_d_in_20_a(array_15_io_d_in_20_a),
    .io_d_in_20_valid_a(array_15_io_d_in_20_valid_a),
    .io_d_in_20_b(array_15_io_d_in_20_b),
    .io_d_in_20_valid_b(array_15_io_d_in_20_valid_b),
    .io_d_in_21_a(array_15_io_d_in_21_a),
    .io_d_in_21_valid_a(array_15_io_d_in_21_valid_a),
    .io_d_in_21_b(array_15_io_d_in_21_b),
    .io_d_in_21_valid_b(array_15_io_d_in_21_valid_b),
    .io_d_in_22_a(array_15_io_d_in_22_a),
    .io_d_in_22_valid_a(array_15_io_d_in_22_valid_a),
    .io_d_in_22_b(array_15_io_d_in_22_b),
    .io_d_in_22_valid_b(array_15_io_d_in_22_valid_b),
    .io_d_in_23_a(array_15_io_d_in_23_a),
    .io_d_in_23_valid_a(array_15_io_d_in_23_valid_a),
    .io_d_in_23_b(array_15_io_d_in_23_b),
    .io_d_in_23_valid_b(array_15_io_d_in_23_valid_b),
    .io_d_in_24_a(array_15_io_d_in_24_a),
    .io_d_in_24_valid_a(array_15_io_d_in_24_valid_a),
    .io_d_in_24_b(array_15_io_d_in_24_b),
    .io_d_in_24_valid_b(array_15_io_d_in_24_valid_b),
    .io_d_in_25_a(array_15_io_d_in_25_a),
    .io_d_in_25_valid_a(array_15_io_d_in_25_valid_a),
    .io_d_in_25_b(array_15_io_d_in_25_b),
    .io_d_in_25_valid_b(array_15_io_d_in_25_valid_b),
    .io_d_in_26_a(array_15_io_d_in_26_a),
    .io_d_in_26_valid_a(array_15_io_d_in_26_valid_a),
    .io_d_in_26_b(array_15_io_d_in_26_b),
    .io_d_in_26_valid_b(array_15_io_d_in_26_valid_b),
    .io_d_in_27_a(array_15_io_d_in_27_a),
    .io_d_in_27_valid_a(array_15_io_d_in_27_valid_a),
    .io_d_in_27_b(array_15_io_d_in_27_b),
    .io_d_in_27_valid_b(array_15_io_d_in_27_valid_b),
    .io_d_in_28_a(array_15_io_d_in_28_a),
    .io_d_in_28_valid_a(array_15_io_d_in_28_valid_a),
    .io_d_in_28_b(array_15_io_d_in_28_b),
    .io_d_in_28_valid_b(array_15_io_d_in_28_valid_b),
    .io_d_in_29_a(array_15_io_d_in_29_a),
    .io_d_in_29_valid_a(array_15_io_d_in_29_valid_a),
    .io_d_in_29_b(array_15_io_d_in_29_b),
    .io_d_in_29_valid_b(array_15_io_d_in_29_valid_b),
    .io_d_in_30_a(array_15_io_d_in_30_a),
    .io_d_in_30_valid_a(array_15_io_d_in_30_valid_a),
    .io_d_in_30_b(array_15_io_d_in_30_b),
    .io_d_in_30_valid_b(array_15_io_d_in_30_valid_b),
    .io_d_in_31_a(array_15_io_d_in_31_a),
    .io_d_in_31_valid_a(array_15_io_d_in_31_valid_a),
    .io_d_in_31_b(array_15_io_d_in_31_b),
    .io_d_in_31_valid_b(array_15_io_d_in_31_valid_b),
    .io_d_out_0_a(array_15_io_d_out_0_a),
    .io_d_out_0_valid_a(array_15_io_d_out_0_valid_a),
    .io_d_out_0_b(array_15_io_d_out_0_b),
    .io_d_out_0_valid_b(array_15_io_d_out_0_valid_b),
    .io_d_out_1_a(array_15_io_d_out_1_a),
    .io_d_out_1_valid_a(array_15_io_d_out_1_valid_a),
    .io_d_out_1_b(array_15_io_d_out_1_b),
    .io_d_out_1_valid_b(array_15_io_d_out_1_valid_b),
    .io_d_out_2_a(array_15_io_d_out_2_a),
    .io_d_out_2_valid_a(array_15_io_d_out_2_valid_a),
    .io_d_out_2_b(array_15_io_d_out_2_b),
    .io_d_out_2_valid_b(array_15_io_d_out_2_valid_b),
    .io_d_out_3_a(array_15_io_d_out_3_a),
    .io_d_out_3_valid_a(array_15_io_d_out_3_valid_a),
    .io_d_out_3_b(array_15_io_d_out_3_b),
    .io_d_out_3_valid_b(array_15_io_d_out_3_valid_b),
    .io_d_out_4_a(array_15_io_d_out_4_a),
    .io_d_out_4_valid_a(array_15_io_d_out_4_valid_a),
    .io_d_out_4_b(array_15_io_d_out_4_b),
    .io_d_out_4_valid_b(array_15_io_d_out_4_valid_b),
    .io_d_out_5_a(array_15_io_d_out_5_a),
    .io_d_out_5_valid_a(array_15_io_d_out_5_valid_a),
    .io_d_out_5_b(array_15_io_d_out_5_b),
    .io_d_out_5_valid_b(array_15_io_d_out_5_valid_b),
    .io_d_out_6_a(array_15_io_d_out_6_a),
    .io_d_out_6_valid_a(array_15_io_d_out_6_valid_a),
    .io_d_out_6_b(array_15_io_d_out_6_b),
    .io_d_out_6_valid_b(array_15_io_d_out_6_valid_b),
    .io_d_out_7_a(array_15_io_d_out_7_a),
    .io_d_out_7_valid_a(array_15_io_d_out_7_valid_a),
    .io_d_out_7_b(array_15_io_d_out_7_b),
    .io_d_out_7_valid_b(array_15_io_d_out_7_valid_b),
    .io_d_out_8_a(array_15_io_d_out_8_a),
    .io_d_out_8_valid_a(array_15_io_d_out_8_valid_a),
    .io_d_out_8_b(array_15_io_d_out_8_b),
    .io_d_out_8_valid_b(array_15_io_d_out_8_valid_b),
    .io_d_out_9_a(array_15_io_d_out_9_a),
    .io_d_out_9_valid_a(array_15_io_d_out_9_valid_a),
    .io_d_out_9_b(array_15_io_d_out_9_b),
    .io_d_out_9_valid_b(array_15_io_d_out_9_valid_b),
    .io_d_out_10_a(array_15_io_d_out_10_a),
    .io_d_out_10_valid_a(array_15_io_d_out_10_valid_a),
    .io_d_out_10_b(array_15_io_d_out_10_b),
    .io_d_out_10_valid_b(array_15_io_d_out_10_valid_b),
    .io_d_out_11_a(array_15_io_d_out_11_a),
    .io_d_out_11_valid_a(array_15_io_d_out_11_valid_a),
    .io_d_out_11_b(array_15_io_d_out_11_b),
    .io_d_out_11_valid_b(array_15_io_d_out_11_valid_b),
    .io_d_out_12_a(array_15_io_d_out_12_a),
    .io_d_out_12_valid_a(array_15_io_d_out_12_valid_a),
    .io_d_out_12_b(array_15_io_d_out_12_b),
    .io_d_out_12_valid_b(array_15_io_d_out_12_valid_b),
    .io_d_out_13_a(array_15_io_d_out_13_a),
    .io_d_out_13_valid_a(array_15_io_d_out_13_valid_a),
    .io_d_out_13_b(array_15_io_d_out_13_b),
    .io_d_out_13_valid_b(array_15_io_d_out_13_valid_b),
    .io_d_out_14_a(array_15_io_d_out_14_a),
    .io_d_out_14_valid_a(array_15_io_d_out_14_valid_a),
    .io_d_out_14_b(array_15_io_d_out_14_b),
    .io_d_out_14_valid_b(array_15_io_d_out_14_valid_b),
    .io_d_out_15_a(array_15_io_d_out_15_a),
    .io_d_out_15_valid_a(array_15_io_d_out_15_valid_a),
    .io_d_out_15_b(array_15_io_d_out_15_b),
    .io_d_out_15_valid_b(array_15_io_d_out_15_valid_b),
    .io_d_out_16_a(array_15_io_d_out_16_a),
    .io_d_out_16_valid_a(array_15_io_d_out_16_valid_a),
    .io_d_out_16_b(array_15_io_d_out_16_b),
    .io_d_out_16_valid_b(array_15_io_d_out_16_valid_b),
    .io_d_out_17_a(array_15_io_d_out_17_a),
    .io_d_out_17_valid_a(array_15_io_d_out_17_valid_a),
    .io_d_out_17_b(array_15_io_d_out_17_b),
    .io_d_out_17_valid_b(array_15_io_d_out_17_valid_b),
    .io_d_out_18_a(array_15_io_d_out_18_a),
    .io_d_out_18_valid_a(array_15_io_d_out_18_valid_a),
    .io_d_out_18_b(array_15_io_d_out_18_b),
    .io_d_out_18_valid_b(array_15_io_d_out_18_valid_b),
    .io_d_out_19_a(array_15_io_d_out_19_a),
    .io_d_out_19_valid_a(array_15_io_d_out_19_valid_a),
    .io_d_out_19_b(array_15_io_d_out_19_b),
    .io_d_out_19_valid_b(array_15_io_d_out_19_valid_b),
    .io_d_out_20_a(array_15_io_d_out_20_a),
    .io_d_out_20_valid_a(array_15_io_d_out_20_valid_a),
    .io_d_out_20_b(array_15_io_d_out_20_b),
    .io_d_out_20_valid_b(array_15_io_d_out_20_valid_b),
    .io_d_out_21_a(array_15_io_d_out_21_a),
    .io_d_out_21_valid_a(array_15_io_d_out_21_valid_a),
    .io_d_out_21_b(array_15_io_d_out_21_b),
    .io_d_out_21_valid_b(array_15_io_d_out_21_valid_b),
    .io_d_out_22_a(array_15_io_d_out_22_a),
    .io_d_out_22_valid_a(array_15_io_d_out_22_valid_a),
    .io_d_out_22_b(array_15_io_d_out_22_b),
    .io_d_out_22_valid_b(array_15_io_d_out_22_valid_b),
    .io_d_out_23_a(array_15_io_d_out_23_a),
    .io_d_out_23_valid_a(array_15_io_d_out_23_valid_a),
    .io_d_out_23_b(array_15_io_d_out_23_b),
    .io_d_out_23_valid_b(array_15_io_d_out_23_valid_b),
    .io_d_out_24_a(array_15_io_d_out_24_a),
    .io_d_out_24_valid_a(array_15_io_d_out_24_valid_a),
    .io_d_out_24_b(array_15_io_d_out_24_b),
    .io_d_out_24_valid_b(array_15_io_d_out_24_valid_b),
    .io_d_out_25_a(array_15_io_d_out_25_a),
    .io_d_out_25_valid_a(array_15_io_d_out_25_valid_a),
    .io_d_out_25_b(array_15_io_d_out_25_b),
    .io_d_out_25_valid_b(array_15_io_d_out_25_valid_b),
    .io_d_out_26_a(array_15_io_d_out_26_a),
    .io_d_out_26_valid_a(array_15_io_d_out_26_valid_a),
    .io_d_out_26_b(array_15_io_d_out_26_b),
    .io_d_out_26_valid_b(array_15_io_d_out_26_valid_b),
    .io_d_out_27_a(array_15_io_d_out_27_a),
    .io_d_out_27_valid_a(array_15_io_d_out_27_valid_a),
    .io_d_out_27_b(array_15_io_d_out_27_b),
    .io_d_out_27_valid_b(array_15_io_d_out_27_valid_b),
    .io_d_out_28_a(array_15_io_d_out_28_a),
    .io_d_out_28_valid_a(array_15_io_d_out_28_valid_a),
    .io_d_out_28_b(array_15_io_d_out_28_b),
    .io_d_out_28_valid_b(array_15_io_d_out_28_valid_b),
    .io_d_out_29_a(array_15_io_d_out_29_a),
    .io_d_out_29_valid_a(array_15_io_d_out_29_valid_a),
    .io_d_out_29_b(array_15_io_d_out_29_b),
    .io_d_out_29_valid_b(array_15_io_d_out_29_valid_b),
    .io_d_out_30_a(array_15_io_d_out_30_a),
    .io_d_out_30_valid_a(array_15_io_d_out_30_valid_a),
    .io_d_out_30_b(array_15_io_d_out_30_b),
    .io_d_out_30_valid_b(array_15_io_d_out_30_valid_b),
    .io_d_out_31_a(array_15_io_d_out_31_a),
    .io_d_out_31_valid_a(array_15_io_d_out_31_valid_a),
    .io_d_out_31_b(array_15_io_d_out_31_b),
    .io_d_out_31_valid_b(array_15_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_15_io_wr_en_mem1),
    .io_wr_en_mem2(array_15_io_wr_en_mem2),
    .io_wr_en_mem3(array_15_io_wr_en_mem3),
    .io_wr_en_mem4(array_15_io_wr_en_mem4),
    .io_wr_en_mem5(array_15_io_wr_en_mem5),
    .io_wr_en_mem6(array_15_io_wr_en_mem6),
    .io_wr_instr_mem1(array_15_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_15_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_15_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_15_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_15_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_15_io_wr_instr_mem6),
    .io_PC1_in(array_15_io_PC1_in),
    .io_PC6_out(array_15_io_PC6_out),
    .io_Addr_in(array_15_io_Addr_in),
    .io_Addr_out(array_15_io_Addr_out)
  );
  BuildingBlockNew array_16 ( // @[BP.scala 45:51]
    .clock(array_16_clock),
    .reset(array_16_reset),
    .io_d_in_0_a(array_16_io_d_in_0_a),
    .io_d_in_0_valid_a(array_16_io_d_in_0_valid_a),
    .io_d_in_0_b(array_16_io_d_in_0_b),
    .io_d_in_0_valid_b(array_16_io_d_in_0_valid_b),
    .io_d_in_1_a(array_16_io_d_in_1_a),
    .io_d_in_1_valid_a(array_16_io_d_in_1_valid_a),
    .io_d_in_1_b(array_16_io_d_in_1_b),
    .io_d_in_1_valid_b(array_16_io_d_in_1_valid_b),
    .io_d_in_2_a(array_16_io_d_in_2_a),
    .io_d_in_2_valid_a(array_16_io_d_in_2_valid_a),
    .io_d_in_2_b(array_16_io_d_in_2_b),
    .io_d_in_2_valid_b(array_16_io_d_in_2_valid_b),
    .io_d_in_3_a(array_16_io_d_in_3_a),
    .io_d_in_3_valid_a(array_16_io_d_in_3_valid_a),
    .io_d_in_3_b(array_16_io_d_in_3_b),
    .io_d_in_3_valid_b(array_16_io_d_in_3_valid_b),
    .io_d_in_4_a(array_16_io_d_in_4_a),
    .io_d_in_4_valid_a(array_16_io_d_in_4_valid_a),
    .io_d_in_4_b(array_16_io_d_in_4_b),
    .io_d_in_4_valid_b(array_16_io_d_in_4_valid_b),
    .io_d_in_5_a(array_16_io_d_in_5_a),
    .io_d_in_5_valid_a(array_16_io_d_in_5_valid_a),
    .io_d_in_5_b(array_16_io_d_in_5_b),
    .io_d_in_5_valid_b(array_16_io_d_in_5_valid_b),
    .io_d_in_6_a(array_16_io_d_in_6_a),
    .io_d_in_6_valid_a(array_16_io_d_in_6_valid_a),
    .io_d_in_6_b(array_16_io_d_in_6_b),
    .io_d_in_6_valid_b(array_16_io_d_in_6_valid_b),
    .io_d_in_7_a(array_16_io_d_in_7_a),
    .io_d_in_7_valid_a(array_16_io_d_in_7_valid_a),
    .io_d_in_7_b(array_16_io_d_in_7_b),
    .io_d_in_7_valid_b(array_16_io_d_in_7_valid_b),
    .io_d_in_8_a(array_16_io_d_in_8_a),
    .io_d_in_8_valid_a(array_16_io_d_in_8_valid_a),
    .io_d_in_8_b(array_16_io_d_in_8_b),
    .io_d_in_8_valid_b(array_16_io_d_in_8_valid_b),
    .io_d_in_9_a(array_16_io_d_in_9_a),
    .io_d_in_9_valid_a(array_16_io_d_in_9_valid_a),
    .io_d_in_9_b(array_16_io_d_in_9_b),
    .io_d_in_9_valid_b(array_16_io_d_in_9_valid_b),
    .io_d_in_10_a(array_16_io_d_in_10_a),
    .io_d_in_10_valid_a(array_16_io_d_in_10_valid_a),
    .io_d_in_10_b(array_16_io_d_in_10_b),
    .io_d_in_10_valid_b(array_16_io_d_in_10_valid_b),
    .io_d_in_11_a(array_16_io_d_in_11_a),
    .io_d_in_11_valid_a(array_16_io_d_in_11_valid_a),
    .io_d_in_11_b(array_16_io_d_in_11_b),
    .io_d_in_11_valid_b(array_16_io_d_in_11_valid_b),
    .io_d_in_12_a(array_16_io_d_in_12_a),
    .io_d_in_12_valid_a(array_16_io_d_in_12_valid_a),
    .io_d_in_12_b(array_16_io_d_in_12_b),
    .io_d_in_12_valid_b(array_16_io_d_in_12_valid_b),
    .io_d_in_13_a(array_16_io_d_in_13_a),
    .io_d_in_13_valid_a(array_16_io_d_in_13_valid_a),
    .io_d_in_13_b(array_16_io_d_in_13_b),
    .io_d_in_13_valid_b(array_16_io_d_in_13_valid_b),
    .io_d_in_14_a(array_16_io_d_in_14_a),
    .io_d_in_14_valid_a(array_16_io_d_in_14_valid_a),
    .io_d_in_14_b(array_16_io_d_in_14_b),
    .io_d_in_14_valid_b(array_16_io_d_in_14_valid_b),
    .io_d_in_15_a(array_16_io_d_in_15_a),
    .io_d_in_15_valid_a(array_16_io_d_in_15_valid_a),
    .io_d_in_15_b(array_16_io_d_in_15_b),
    .io_d_in_15_valid_b(array_16_io_d_in_15_valid_b),
    .io_d_in_16_a(array_16_io_d_in_16_a),
    .io_d_in_16_valid_a(array_16_io_d_in_16_valid_a),
    .io_d_in_16_b(array_16_io_d_in_16_b),
    .io_d_in_16_valid_b(array_16_io_d_in_16_valid_b),
    .io_d_in_17_a(array_16_io_d_in_17_a),
    .io_d_in_17_valid_a(array_16_io_d_in_17_valid_a),
    .io_d_in_17_b(array_16_io_d_in_17_b),
    .io_d_in_17_valid_b(array_16_io_d_in_17_valid_b),
    .io_d_in_18_a(array_16_io_d_in_18_a),
    .io_d_in_18_valid_a(array_16_io_d_in_18_valid_a),
    .io_d_in_18_b(array_16_io_d_in_18_b),
    .io_d_in_18_valid_b(array_16_io_d_in_18_valid_b),
    .io_d_in_19_a(array_16_io_d_in_19_a),
    .io_d_in_19_valid_a(array_16_io_d_in_19_valid_a),
    .io_d_in_19_b(array_16_io_d_in_19_b),
    .io_d_in_19_valid_b(array_16_io_d_in_19_valid_b),
    .io_d_in_20_a(array_16_io_d_in_20_a),
    .io_d_in_20_valid_a(array_16_io_d_in_20_valid_a),
    .io_d_in_20_b(array_16_io_d_in_20_b),
    .io_d_in_20_valid_b(array_16_io_d_in_20_valid_b),
    .io_d_in_21_a(array_16_io_d_in_21_a),
    .io_d_in_21_valid_a(array_16_io_d_in_21_valid_a),
    .io_d_in_21_b(array_16_io_d_in_21_b),
    .io_d_in_21_valid_b(array_16_io_d_in_21_valid_b),
    .io_d_in_22_a(array_16_io_d_in_22_a),
    .io_d_in_22_valid_a(array_16_io_d_in_22_valid_a),
    .io_d_in_22_b(array_16_io_d_in_22_b),
    .io_d_in_22_valid_b(array_16_io_d_in_22_valid_b),
    .io_d_in_23_a(array_16_io_d_in_23_a),
    .io_d_in_23_valid_a(array_16_io_d_in_23_valid_a),
    .io_d_in_23_b(array_16_io_d_in_23_b),
    .io_d_in_23_valid_b(array_16_io_d_in_23_valid_b),
    .io_d_in_24_a(array_16_io_d_in_24_a),
    .io_d_in_24_valid_a(array_16_io_d_in_24_valid_a),
    .io_d_in_24_b(array_16_io_d_in_24_b),
    .io_d_in_24_valid_b(array_16_io_d_in_24_valid_b),
    .io_d_in_25_a(array_16_io_d_in_25_a),
    .io_d_in_25_valid_a(array_16_io_d_in_25_valid_a),
    .io_d_in_25_b(array_16_io_d_in_25_b),
    .io_d_in_25_valid_b(array_16_io_d_in_25_valid_b),
    .io_d_in_26_a(array_16_io_d_in_26_a),
    .io_d_in_26_valid_a(array_16_io_d_in_26_valid_a),
    .io_d_in_26_b(array_16_io_d_in_26_b),
    .io_d_in_26_valid_b(array_16_io_d_in_26_valid_b),
    .io_d_in_27_a(array_16_io_d_in_27_a),
    .io_d_in_27_valid_a(array_16_io_d_in_27_valid_a),
    .io_d_in_27_b(array_16_io_d_in_27_b),
    .io_d_in_27_valid_b(array_16_io_d_in_27_valid_b),
    .io_d_in_28_a(array_16_io_d_in_28_a),
    .io_d_in_28_valid_a(array_16_io_d_in_28_valid_a),
    .io_d_in_28_b(array_16_io_d_in_28_b),
    .io_d_in_28_valid_b(array_16_io_d_in_28_valid_b),
    .io_d_in_29_a(array_16_io_d_in_29_a),
    .io_d_in_29_valid_a(array_16_io_d_in_29_valid_a),
    .io_d_in_29_b(array_16_io_d_in_29_b),
    .io_d_in_29_valid_b(array_16_io_d_in_29_valid_b),
    .io_d_in_30_a(array_16_io_d_in_30_a),
    .io_d_in_30_valid_a(array_16_io_d_in_30_valid_a),
    .io_d_in_30_b(array_16_io_d_in_30_b),
    .io_d_in_30_valid_b(array_16_io_d_in_30_valid_b),
    .io_d_in_31_a(array_16_io_d_in_31_a),
    .io_d_in_31_valid_a(array_16_io_d_in_31_valid_a),
    .io_d_in_31_b(array_16_io_d_in_31_b),
    .io_d_in_31_valid_b(array_16_io_d_in_31_valid_b),
    .io_d_out_0_a(array_16_io_d_out_0_a),
    .io_d_out_0_valid_a(array_16_io_d_out_0_valid_a),
    .io_d_out_0_b(array_16_io_d_out_0_b),
    .io_d_out_0_valid_b(array_16_io_d_out_0_valid_b),
    .io_d_out_1_a(array_16_io_d_out_1_a),
    .io_d_out_1_valid_a(array_16_io_d_out_1_valid_a),
    .io_d_out_1_b(array_16_io_d_out_1_b),
    .io_d_out_1_valid_b(array_16_io_d_out_1_valid_b),
    .io_d_out_2_a(array_16_io_d_out_2_a),
    .io_d_out_2_valid_a(array_16_io_d_out_2_valid_a),
    .io_d_out_2_b(array_16_io_d_out_2_b),
    .io_d_out_2_valid_b(array_16_io_d_out_2_valid_b),
    .io_d_out_3_a(array_16_io_d_out_3_a),
    .io_d_out_3_valid_a(array_16_io_d_out_3_valid_a),
    .io_d_out_3_b(array_16_io_d_out_3_b),
    .io_d_out_3_valid_b(array_16_io_d_out_3_valid_b),
    .io_d_out_4_a(array_16_io_d_out_4_a),
    .io_d_out_4_valid_a(array_16_io_d_out_4_valid_a),
    .io_d_out_4_b(array_16_io_d_out_4_b),
    .io_d_out_4_valid_b(array_16_io_d_out_4_valid_b),
    .io_d_out_5_a(array_16_io_d_out_5_a),
    .io_d_out_5_valid_a(array_16_io_d_out_5_valid_a),
    .io_d_out_5_b(array_16_io_d_out_5_b),
    .io_d_out_5_valid_b(array_16_io_d_out_5_valid_b),
    .io_d_out_6_a(array_16_io_d_out_6_a),
    .io_d_out_6_valid_a(array_16_io_d_out_6_valid_a),
    .io_d_out_6_b(array_16_io_d_out_6_b),
    .io_d_out_6_valid_b(array_16_io_d_out_6_valid_b),
    .io_d_out_7_a(array_16_io_d_out_7_a),
    .io_d_out_7_valid_a(array_16_io_d_out_7_valid_a),
    .io_d_out_7_b(array_16_io_d_out_7_b),
    .io_d_out_7_valid_b(array_16_io_d_out_7_valid_b),
    .io_d_out_8_a(array_16_io_d_out_8_a),
    .io_d_out_8_valid_a(array_16_io_d_out_8_valid_a),
    .io_d_out_8_b(array_16_io_d_out_8_b),
    .io_d_out_8_valid_b(array_16_io_d_out_8_valid_b),
    .io_d_out_9_a(array_16_io_d_out_9_a),
    .io_d_out_9_valid_a(array_16_io_d_out_9_valid_a),
    .io_d_out_9_b(array_16_io_d_out_9_b),
    .io_d_out_9_valid_b(array_16_io_d_out_9_valid_b),
    .io_d_out_10_a(array_16_io_d_out_10_a),
    .io_d_out_10_valid_a(array_16_io_d_out_10_valid_a),
    .io_d_out_10_b(array_16_io_d_out_10_b),
    .io_d_out_10_valid_b(array_16_io_d_out_10_valid_b),
    .io_d_out_11_a(array_16_io_d_out_11_a),
    .io_d_out_11_valid_a(array_16_io_d_out_11_valid_a),
    .io_d_out_11_b(array_16_io_d_out_11_b),
    .io_d_out_11_valid_b(array_16_io_d_out_11_valid_b),
    .io_d_out_12_a(array_16_io_d_out_12_a),
    .io_d_out_12_valid_a(array_16_io_d_out_12_valid_a),
    .io_d_out_12_b(array_16_io_d_out_12_b),
    .io_d_out_12_valid_b(array_16_io_d_out_12_valid_b),
    .io_d_out_13_a(array_16_io_d_out_13_a),
    .io_d_out_13_valid_a(array_16_io_d_out_13_valid_a),
    .io_d_out_13_b(array_16_io_d_out_13_b),
    .io_d_out_13_valid_b(array_16_io_d_out_13_valid_b),
    .io_d_out_14_a(array_16_io_d_out_14_a),
    .io_d_out_14_valid_a(array_16_io_d_out_14_valid_a),
    .io_d_out_14_b(array_16_io_d_out_14_b),
    .io_d_out_14_valid_b(array_16_io_d_out_14_valid_b),
    .io_d_out_15_a(array_16_io_d_out_15_a),
    .io_d_out_15_valid_a(array_16_io_d_out_15_valid_a),
    .io_d_out_15_b(array_16_io_d_out_15_b),
    .io_d_out_15_valid_b(array_16_io_d_out_15_valid_b),
    .io_d_out_16_a(array_16_io_d_out_16_a),
    .io_d_out_16_valid_a(array_16_io_d_out_16_valid_a),
    .io_d_out_16_b(array_16_io_d_out_16_b),
    .io_d_out_16_valid_b(array_16_io_d_out_16_valid_b),
    .io_d_out_17_a(array_16_io_d_out_17_a),
    .io_d_out_17_valid_a(array_16_io_d_out_17_valid_a),
    .io_d_out_17_b(array_16_io_d_out_17_b),
    .io_d_out_17_valid_b(array_16_io_d_out_17_valid_b),
    .io_d_out_18_a(array_16_io_d_out_18_a),
    .io_d_out_18_valid_a(array_16_io_d_out_18_valid_a),
    .io_d_out_18_b(array_16_io_d_out_18_b),
    .io_d_out_18_valid_b(array_16_io_d_out_18_valid_b),
    .io_d_out_19_a(array_16_io_d_out_19_a),
    .io_d_out_19_valid_a(array_16_io_d_out_19_valid_a),
    .io_d_out_19_b(array_16_io_d_out_19_b),
    .io_d_out_19_valid_b(array_16_io_d_out_19_valid_b),
    .io_d_out_20_a(array_16_io_d_out_20_a),
    .io_d_out_20_valid_a(array_16_io_d_out_20_valid_a),
    .io_d_out_20_b(array_16_io_d_out_20_b),
    .io_d_out_20_valid_b(array_16_io_d_out_20_valid_b),
    .io_d_out_21_a(array_16_io_d_out_21_a),
    .io_d_out_21_valid_a(array_16_io_d_out_21_valid_a),
    .io_d_out_21_b(array_16_io_d_out_21_b),
    .io_d_out_21_valid_b(array_16_io_d_out_21_valid_b),
    .io_d_out_22_a(array_16_io_d_out_22_a),
    .io_d_out_22_valid_a(array_16_io_d_out_22_valid_a),
    .io_d_out_22_b(array_16_io_d_out_22_b),
    .io_d_out_22_valid_b(array_16_io_d_out_22_valid_b),
    .io_d_out_23_a(array_16_io_d_out_23_a),
    .io_d_out_23_valid_a(array_16_io_d_out_23_valid_a),
    .io_d_out_23_b(array_16_io_d_out_23_b),
    .io_d_out_23_valid_b(array_16_io_d_out_23_valid_b),
    .io_d_out_24_a(array_16_io_d_out_24_a),
    .io_d_out_24_valid_a(array_16_io_d_out_24_valid_a),
    .io_d_out_24_b(array_16_io_d_out_24_b),
    .io_d_out_24_valid_b(array_16_io_d_out_24_valid_b),
    .io_d_out_25_a(array_16_io_d_out_25_a),
    .io_d_out_25_valid_a(array_16_io_d_out_25_valid_a),
    .io_d_out_25_b(array_16_io_d_out_25_b),
    .io_d_out_25_valid_b(array_16_io_d_out_25_valid_b),
    .io_d_out_26_a(array_16_io_d_out_26_a),
    .io_d_out_26_valid_a(array_16_io_d_out_26_valid_a),
    .io_d_out_26_b(array_16_io_d_out_26_b),
    .io_d_out_26_valid_b(array_16_io_d_out_26_valid_b),
    .io_d_out_27_a(array_16_io_d_out_27_a),
    .io_d_out_27_valid_a(array_16_io_d_out_27_valid_a),
    .io_d_out_27_b(array_16_io_d_out_27_b),
    .io_d_out_27_valid_b(array_16_io_d_out_27_valid_b),
    .io_d_out_28_a(array_16_io_d_out_28_a),
    .io_d_out_28_valid_a(array_16_io_d_out_28_valid_a),
    .io_d_out_28_b(array_16_io_d_out_28_b),
    .io_d_out_28_valid_b(array_16_io_d_out_28_valid_b),
    .io_d_out_29_a(array_16_io_d_out_29_a),
    .io_d_out_29_valid_a(array_16_io_d_out_29_valid_a),
    .io_d_out_29_b(array_16_io_d_out_29_b),
    .io_d_out_29_valid_b(array_16_io_d_out_29_valid_b),
    .io_d_out_30_a(array_16_io_d_out_30_a),
    .io_d_out_30_valid_a(array_16_io_d_out_30_valid_a),
    .io_d_out_30_b(array_16_io_d_out_30_b),
    .io_d_out_30_valid_b(array_16_io_d_out_30_valid_b),
    .io_d_out_31_a(array_16_io_d_out_31_a),
    .io_d_out_31_valid_a(array_16_io_d_out_31_valid_a),
    .io_d_out_31_b(array_16_io_d_out_31_b),
    .io_d_out_31_valid_b(array_16_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_16_io_wr_en_mem1),
    .io_wr_en_mem2(array_16_io_wr_en_mem2),
    .io_wr_en_mem3(array_16_io_wr_en_mem3),
    .io_wr_en_mem4(array_16_io_wr_en_mem4),
    .io_wr_en_mem5(array_16_io_wr_en_mem5),
    .io_wr_en_mem6(array_16_io_wr_en_mem6),
    .io_wr_instr_mem1(array_16_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_16_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_16_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_16_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_16_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_16_io_wr_instr_mem6),
    .io_PC1_in(array_16_io_PC1_in),
    .io_PC6_out(array_16_io_PC6_out),
    .io_Addr_in(array_16_io_Addr_in),
    .io_Addr_out(array_16_io_Addr_out)
  );
  BuildingBlockNew array_17 ( // @[BP.scala 45:51]
    .clock(array_17_clock),
    .reset(array_17_reset),
    .io_d_in_0_a(array_17_io_d_in_0_a),
    .io_d_in_0_valid_a(array_17_io_d_in_0_valid_a),
    .io_d_in_0_b(array_17_io_d_in_0_b),
    .io_d_in_0_valid_b(array_17_io_d_in_0_valid_b),
    .io_d_in_1_a(array_17_io_d_in_1_a),
    .io_d_in_1_valid_a(array_17_io_d_in_1_valid_a),
    .io_d_in_1_b(array_17_io_d_in_1_b),
    .io_d_in_1_valid_b(array_17_io_d_in_1_valid_b),
    .io_d_in_2_a(array_17_io_d_in_2_a),
    .io_d_in_2_valid_a(array_17_io_d_in_2_valid_a),
    .io_d_in_2_b(array_17_io_d_in_2_b),
    .io_d_in_2_valid_b(array_17_io_d_in_2_valid_b),
    .io_d_in_3_a(array_17_io_d_in_3_a),
    .io_d_in_3_valid_a(array_17_io_d_in_3_valid_a),
    .io_d_in_3_b(array_17_io_d_in_3_b),
    .io_d_in_3_valid_b(array_17_io_d_in_3_valid_b),
    .io_d_in_4_a(array_17_io_d_in_4_a),
    .io_d_in_4_valid_a(array_17_io_d_in_4_valid_a),
    .io_d_in_4_b(array_17_io_d_in_4_b),
    .io_d_in_4_valid_b(array_17_io_d_in_4_valid_b),
    .io_d_in_5_a(array_17_io_d_in_5_a),
    .io_d_in_5_valid_a(array_17_io_d_in_5_valid_a),
    .io_d_in_5_b(array_17_io_d_in_5_b),
    .io_d_in_5_valid_b(array_17_io_d_in_5_valid_b),
    .io_d_in_6_a(array_17_io_d_in_6_a),
    .io_d_in_6_valid_a(array_17_io_d_in_6_valid_a),
    .io_d_in_6_b(array_17_io_d_in_6_b),
    .io_d_in_6_valid_b(array_17_io_d_in_6_valid_b),
    .io_d_in_7_a(array_17_io_d_in_7_a),
    .io_d_in_7_valid_a(array_17_io_d_in_7_valid_a),
    .io_d_in_7_b(array_17_io_d_in_7_b),
    .io_d_in_7_valid_b(array_17_io_d_in_7_valid_b),
    .io_d_in_8_a(array_17_io_d_in_8_a),
    .io_d_in_8_valid_a(array_17_io_d_in_8_valid_a),
    .io_d_in_8_b(array_17_io_d_in_8_b),
    .io_d_in_8_valid_b(array_17_io_d_in_8_valid_b),
    .io_d_in_9_a(array_17_io_d_in_9_a),
    .io_d_in_9_valid_a(array_17_io_d_in_9_valid_a),
    .io_d_in_9_b(array_17_io_d_in_9_b),
    .io_d_in_9_valid_b(array_17_io_d_in_9_valid_b),
    .io_d_in_10_a(array_17_io_d_in_10_a),
    .io_d_in_10_valid_a(array_17_io_d_in_10_valid_a),
    .io_d_in_10_b(array_17_io_d_in_10_b),
    .io_d_in_10_valid_b(array_17_io_d_in_10_valid_b),
    .io_d_in_11_a(array_17_io_d_in_11_a),
    .io_d_in_11_valid_a(array_17_io_d_in_11_valid_a),
    .io_d_in_11_b(array_17_io_d_in_11_b),
    .io_d_in_11_valid_b(array_17_io_d_in_11_valid_b),
    .io_d_in_12_a(array_17_io_d_in_12_a),
    .io_d_in_12_valid_a(array_17_io_d_in_12_valid_a),
    .io_d_in_12_b(array_17_io_d_in_12_b),
    .io_d_in_12_valid_b(array_17_io_d_in_12_valid_b),
    .io_d_in_13_a(array_17_io_d_in_13_a),
    .io_d_in_13_valid_a(array_17_io_d_in_13_valid_a),
    .io_d_in_13_b(array_17_io_d_in_13_b),
    .io_d_in_13_valid_b(array_17_io_d_in_13_valid_b),
    .io_d_in_14_a(array_17_io_d_in_14_a),
    .io_d_in_14_valid_a(array_17_io_d_in_14_valid_a),
    .io_d_in_14_b(array_17_io_d_in_14_b),
    .io_d_in_14_valid_b(array_17_io_d_in_14_valid_b),
    .io_d_in_15_a(array_17_io_d_in_15_a),
    .io_d_in_15_valid_a(array_17_io_d_in_15_valid_a),
    .io_d_in_15_b(array_17_io_d_in_15_b),
    .io_d_in_15_valid_b(array_17_io_d_in_15_valid_b),
    .io_d_in_16_a(array_17_io_d_in_16_a),
    .io_d_in_16_valid_a(array_17_io_d_in_16_valid_a),
    .io_d_in_16_b(array_17_io_d_in_16_b),
    .io_d_in_16_valid_b(array_17_io_d_in_16_valid_b),
    .io_d_in_17_a(array_17_io_d_in_17_a),
    .io_d_in_17_valid_a(array_17_io_d_in_17_valid_a),
    .io_d_in_17_b(array_17_io_d_in_17_b),
    .io_d_in_17_valid_b(array_17_io_d_in_17_valid_b),
    .io_d_in_18_a(array_17_io_d_in_18_a),
    .io_d_in_18_valid_a(array_17_io_d_in_18_valid_a),
    .io_d_in_18_b(array_17_io_d_in_18_b),
    .io_d_in_18_valid_b(array_17_io_d_in_18_valid_b),
    .io_d_in_19_a(array_17_io_d_in_19_a),
    .io_d_in_19_valid_a(array_17_io_d_in_19_valid_a),
    .io_d_in_19_b(array_17_io_d_in_19_b),
    .io_d_in_19_valid_b(array_17_io_d_in_19_valid_b),
    .io_d_in_20_a(array_17_io_d_in_20_a),
    .io_d_in_20_valid_a(array_17_io_d_in_20_valid_a),
    .io_d_in_20_b(array_17_io_d_in_20_b),
    .io_d_in_20_valid_b(array_17_io_d_in_20_valid_b),
    .io_d_in_21_a(array_17_io_d_in_21_a),
    .io_d_in_21_valid_a(array_17_io_d_in_21_valid_a),
    .io_d_in_21_b(array_17_io_d_in_21_b),
    .io_d_in_21_valid_b(array_17_io_d_in_21_valid_b),
    .io_d_in_22_a(array_17_io_d_in_22_a),
    .io_d_in_22_valid_a(array_17_io_d_in_22_valid_a),
    .io_d_in_22_b(array_17_io_d_in_22_b),
    .io_d_in_22_valid_b(array_17_io_d_in_22_valid_b),
    .io_d_in_23_a(array_17_io_d_in_23_a),
    .io_d_in_23_valid_a(array_17_io_d_in_23_valid_a),
    .io_d_in_23_b(array_17_io_d_in_23_b),
    .io_d_in_23_valid_b(array_17_io_d_in_23_valid_b),
    .io_d_in_24_a(array_17_io_d_in_24_a),
    .io_d_in_24_valid_a(array_17_io_d_in_24_valid_a),
    .io_d_in_24_b(array_17_io_d_in_24_b),
    .io_d_in_24_valid_b(array_17_io_d_in_24_valid_b),
    .io_d_in_25_a(array_17_io_d_in_25_a),
    .io_d_in_25_valid_a(array_17_io_d_in_25_valid_a),
    .io_d_in_25_b(array_17_io_d_in_25_b),
    .io_d_in_25_valid_b(array_17_io_d_in_25_valid_b),
    .io_d_in_26_a(array_17_io_d_in_26_a),
    .io_d_in_26_valid_a(array_17_io_d_in_26_valid_a),
    .io_d_in_26_b(array_17_io_d_in_26_b),
    .io_d_in_26_valid_b(array_17_io_d_in_26_valid_b),
    .io_d_in_27_a(array_17_io_d_in_27_a),
    .io_d_in_27_valid_a(array_17_io_d_in_27_valid_a),
    .io_d_in_27_b(array_17_io_d_in_27_b),
    .io_d_in_27_valid_b(array_17_io_d_in_27_valid_b),
    .io_d_in_28_a(array_17_io_d_in_28_a),
    .io_d_in_28_valid_a(array_17_io_d_in_28_valid_a),
    .io_d_in_28_b(array_17_io_d_in_28_b),
    .io_d_in_28_valid_b(array_17_io_d_in_28_valid_b),
    .io_d_in_29_a(array_17_io_d_in_29_a),
    .io_d_in_29_valid_a(array_17_io_d_in_29_valid_a),
    .io_d_in_29_b(array_17_io_d_in_29_b),
    .io_d_in_29_valid_b(array_17_io_d_in_29_valid_b),
    .io_d_in_30_a(array_17_io_d_in_30_a),
    .io_d_in_30_valid_a(array_17_io_d_in_30_valid_a),
    .io_d_in_30_b(array_17_io_d_in_30_b),
    .io_d_in_30_valid_b(array_17_io_d_in_30_valid_b),
    .io_d_in_31_a(array_17_io_d_in_31_a),
    .io_d_in_31_valid_a(array_17_io_d_in_31_valid_a),
    .io_d_in_31_b(array_17_io_d_in_31_b),
    .io_d_in_31_valid_b(array_17_io_d_in_31_valid_b),
    .io_d_out_0_a(array_17_io_d_out_0_a),
    .io_d_out_0_valid_a(array_17_io_d_out_0_valid_a),
    .io_d_out_0_b(array_17_io_d_out_0_b),
    .io_d_out_0_valid_b(array_17_io_d_out_0_valid_b),
    .io_d_out_1_a(array_17_io_d_out_1_a),
    .io_d_out_1_valid_a(array_17_io_d_out_1_valid_a),
    .io_d_out_1_b(array_17_io_d_out_1_b),
    .io_d_out_1_valid_b(array_17_io_d_out_1_valid_b),
    .io_d_out_2_a(array_17_io_d_out_2_a),
    .io_d_out_2_valid_a(array_17_io_d_out_2_valid_a),
    .io_d_out_2_b(array_17_io_d_out_2_b),
    .io_d_out_2_valid_b(array_17_io_d_out_2_valid_b),
    .io_d_out_3_a(array_17_io_d_out_3_a),
    .io_d_out_3_valid_a(array_17_io_d_out_3_valid_a),
    .io_d_out_3_b(array_17_io_d_out_3_b),
    .io_d_out_3_valid_b(array_17_io_d_out_3_valid_b),
    .io_d_out_4_a(array_17_io_d_out_4_a),
    .io_d_out_4_valid_a(array_17_io_d_out_4_valid_a),
    .io_d_out_4_b(array_17_io_d_out_4_b),
    .io_d_out_4_valid_b(array_17_io_d_out_4_valid_b),
    .io_d_out_5_a(array_17_io_d_out_5_a),
    .io_d_out_5_valid_a(array_17_io_d_out_5_valid_a),
    .io_d_out_5_b(array_17_io_d_out_5_b),
    .io_d_out_5_valid_b(array_17_io_d_out_5_valid_b),
    .io_d_out_6_a(array_17_io_d_out_6_a),
    .io_d_out_6_valid_a(array_17_io_d_out_6_valid_a),
    .io_d_out_6_b(array_17_io_d_out_6_b),
    .io_d_out_6_valid_b(array_17_io_d_out_6_valid_b),
    .io_d_out_7_a(array_17_io_d_out_7_a),
    .io_d_out_7_valid_a(array_17_io_d_out_7_valid_a),
    .io_d_out_7_b(array_17_io_d_out_7_b),
    .io_d_out_7_valid_b(array_17_io_d_out_7_valid_b),
    .io_d_out_8_a(array_17_io_d_out_8_a),
    .io_d_out_8_valid_a(array_17_io_d_out_8_valid_a),
    .io_d_out_8_b(array_17_io_d_out_8_b),
    .io_d_out_8_valid_b(array_17_io_d_out_8_valid_b),
    .io_d_out_9_a(array_17_io_d_out_9_a),
    .io_d_out_9_valid_a(array_17_io_d_out_9_valid_a),
    .io_d_out_9_b(array_17_io_d_out_9_b),
    .io_d_out_9_valid_b(array_17_io_d_out_9_valid_b),
    .io_d_out_10_a(array_17_io_d_out_10_a),
    .io_d_out_10_valid_a(array_17_io_d_out_10_valid_a),
    .io_d_out_10_b(array_17_io_d_out_10_b),
    .io_d_out_10_valid_b(array_17_io_d_out_10_valid_b),
    .io_d_out_11_a(array_17_io_d_out_11_a),
    .io_d_out_11_valid_a(array_17_io_d_out_11_valid_a),
    .io_d_out_11_b(array_17_io_d_out_11_b),
    .io_d_out_11_valid_b(array_17_io_d_out_11_valid_b),
    .io_d_out_12_a(array_17_io_d_out_12_a),
    .io_d_out_12_valid_a(array_17_io_d_out_12_valid_a),
    .io_d_out_12_b(array_17_io_d_out_12_b),
    .io_d_out_12_valid_b(array_17_io_d_out_12_valid_b),
    .io_d_out_13_a(array_17_io_d_out_13_a),
    .io_d_out_13_valid_a(array_17_io_d_out_13_valid_a),
    .io_d_out_13_b(array_17_io_d_out_13_b),
    .io_d_out_13_valid_b(array_17_io_d_out_13_valid_b),
    .io_d_out_14_a(array_17_io_d_out_14_a),
    .io_d_out_14_valid_a(array_17_io_d_out_14_valid_a),
    .io_d_out_14_b(array_17_io_d_out_14_b),
    .io_d_out_14_valid_b(array_17_io_d_out_14_valid_b),
    .io_d_out_15_a(array_17_io_d_out_15_a),
    .io_d_out_15_valid_a(array_17_io_d_out_15_valid_a),
    .io_d_out_15_b(array_17_io_d_out_15_b),
    .io_d_out_15_valid_b(array_17_io_d_out_15_valid_b),
    .io_d_out_16_a(array_17_io_d_out_16_a),
    .io_d_out_16_valid_a(array_17_io_d_out_16_valid_a),
    .io_d_out_16_b(array_17_io_d_out_16_b),
    .io_d_out_16_valid_b(array_17_io_d_out_16_valid_b),
    .io_d_out_17_a(array_17_io_d_out_17_a),
    .io_d_out_17_valid_a(array_17_io_d_out_17_valid_a),
    .io_d_out_17_b(array_17_io_d_out_17_b),
    .io_d_out_17_valid_b(array_17_io_d_out_17_valid_b),
    .io_d_out_18_a(array_17_io_d_out_18_a),
    .io_d_out_18_valid_a(array_17_io_d_out_18_valid_a),
    .io_d_out_18_b(array_17_io_d_out_18_b),
    .io_d_out_18_valid_b(array_17_io_d_out_18_valid_b),
    .io_d_out_19_a(array_17_io_d_out_19_a),
    .io_d_out_19_valid_a(array_17_io_d_out_19_valid_a),
    .io_d_out_19_b(array_17_io_d_out_19_b),
    .io_d_out_19_valid_b(array_17_io_d_out_19_valid_b),
    .io_d_out_20_a(array_17_io_d_out_20_a),
    .io_d_out_20_valid_a(array_17_io_d_out_20_valid_a),
    .io_d_out_20_b(array_17_io_d_out_20_b),
    .io_d_out_20_valid_b(array_17_io_d_out_20_valid_b),
    .io_d_out_21_a(array_17_io_d_out_21_a),
    .io_d_out_21_valid_a(array_17_io_d_out_21_valid_a),
    .io_d_out_21_b(array_17_io_d_out_21_b),
    .io_d_out_21_valid_b(array_17_io_d_out_21_valid_b),
    .io_d_out_22_a(array_17_io_d_out_22_a),
    .io_d_out_22_valid_a(array_17_io_d_out_22_valid_a),
    .io_d_out_22_b(array_17_io_d_out_22_b),
    .io_d_out_22_valid_b(array_17_io_d_out_22_valid_b),
    .io_d_out_23_a(array_17_io_d_out_23_a),
    .io_d_out_23_valid_a(array_17_io_d_out_23_valid_a),
    .io_d_out_23_b(array_17_io_d_out_23_b),
    .io_d_out_23_valid_b(array_17_io_d_out_23_valid_b),
    .io_d_out_24_a(array_17_io_d_out_24_a),
    .io_d_out_24_valid_a(array_17_io_d_out_24_valid_a),
    .io_d_out_24_b(array_17_io_d_out_24_b),
    .io_d_out_24_valid_b(array_17_io_d_out_24_valid_b),
    .io_d_out_25_a(array_17_io_d_out_25_a),
    .io_d_out_25_valid_a(array_17_io_d_out_25_valid_a),
    .io_d_out_25_b(array_17_io_d_out_25_b),
    .io_d_out_25_valid_b(array_17_io_d_out_25_valid_b),
    .io_d_out_26_a(array_17_io_d_out_26_a),
    .io_d_out_26_valid_a(array_17_io_d_out_26_valid_a),
    .io_d_out_26_b(array_17_io_d_out_26_b),
    .io_d_out_26_valid_b(array_17_io_d_out_26_valid_b),
    .io_d_out_27_a(array_17_io_d_out_27_a),
    .io_d_out_27_valid_a(array_17_io_d_out_27_valid_a),
    .io_d_out_27_b(array_17_io_d_out_27_b),
    .io_d_out_27_valid_b(array_17_io_d_out_27_valid_b),
    .io_d_out_28_a(array_17_io_d_out_28_a),
    .io_d_out_28_valid_a(array_17_io_d_out_28_valid_a),
    .io_d_out_28_b(array_17_io_d_out_28_b),
    .io_d_out_28_valid_b(array_17_io_d_out_28_valid_b),
    .io_d_out_29_a(array_17_io_d_out_29_a),
    .io_d_out_29_valid_a(array_17_io_d_out_29_valid_a),
    .io_d_out_29_b(array_17_io_d_out_29_b),
    .io_d_out_29_valid_b(array_17_io_d_out_29_valid_b),
    .io_d_out_30_a(array_17_io_d_out_30_a),
    .io_d_out_30_valid_a(array_17_io_d_out_30_valid_a),
    .io_d_out_30_b(array_17_io_d_out_30_b),
    .io_d_out_30_valid_b(array_17_io_d_out_30_valid_b),
    .io_d_out_31_a(array_17_io_d_out_31_a),
    .io_d_out_31_valid_a(array_17_io_d_out_31_valid_a),
    .io_d_out_31_b(array_17_io_d_out_31_b),
    .io_d_out_31_valid_b(array_17_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_17_io_wr_en_mem1),
    .io_wr_en_mem2(array_17_io_wr_en_mem2),
    .io_wr_en_mem3(array_17_io_wr_en_mem3),
    .io_wr_en_mem4(array_17_io_wr_en_mem4),
    .io_wr_en_mem5(array_17_io_wr_en_mem5),
    .io_wr_en_mem6(array_17_io_wr_en_mem6),
    .io_wr_instr_mem1(array_17_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_17_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_17_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_17_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_17_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_17_io_wr_instr_mem6),
    .io_PC1_in(array_17_io_PC1_in),
    .io_PC6_out(array_17_io_PC6_out),
    .io_Addr_in(array_17_io_Addr_in),
    .io_Addr_out(array_17_io_Addr_out)
  );
  BuildingBlockNew array_18 ( // @[BP.scala 45:51]
    .clock(array_18_clock),
    .reset(array_18_reset),
    .io_d_in_0_a(array_18_io_d_in_0_a),
    .io_d_in_0_valid_a(array_18_io_d_in_0_valid_a),
    .io_d_in_0_b(array_18_io_d_in_0_b),
    .io_d_in_0_valid_b(array_18_io_d_in_0_valid_b),
    .io_d_in_1_a(array_18_io_d_in_1_a),
    .io_d_in_1_valid_a(array_18_io_d_in_1_valid_a),
    .io_d_in_1_b(array_18_io_d_in_1_b),
    .io_d_in_1_valid_b(array_18_io_d_in_1_valid_b),
    .io_d_in_2_a(array_18_io_d_in_2_a),
    .io_d_in_2_valid_a(array_18_io_d_in_2_valid_a),
    .io_d_in_2_b(array_18_io_d_in_2_b),
    .io_d_in_2_valid_b(array_18_io_d_in_2_valid_b),
    .io_d_in_3_a(array_18_io_d_in_3_a),
    .io_d_in_3_valid_a(array_18_io_d_in_3_valid_a),
    .io_d_in_3_b(array_18_io_d_in_3_b),
    .io_d_in_3_valid_b(array_18_io_d_in_3_valid_b),
    .io_d_in_4_a(array_18_io_d_in_4_a),
    .io_d_in_4_valid_a(array_18_io_d_in_4_valid_a),
    .io_d_in_4_b(array_18_io_d_in_4_b),
    .io_d_in_4_valid_b(array_18_io_d_in_4_valid_b),
    .io_d_in_5_a(array_18_io_d_in_5_a),
    .io_d_in_5_valid_a(array_18_io_d_in_5_valid_a),
    .io_d_in_5_b(array_18_io_d_in_5_b),
    .io_d_in_5_valid_b(array_18_io_d_in_5_valid_b),
    .io_d_in_6_a(array_18_io_d_in_6_a),
    .io_d_in_6_valid_a(array_18_io_d_in_6_valid_a),
    .io_d_in_6_b(array_18_io_d_in_6_b),
    .io_d_in_6_valid_b(array_18_io_d_in_6_valid_b),
    .io_d_in_7_a(array_18_io_d_in_7_a),
    .io_d_in_7_valid_a(array_18_io_d_in_7_valid_a),
    .io_d_in_7_b(array_18_io_d_in_7_b),
    .io_d_in_7_valid_b(array_18_io_d_in_7_valid_b),
    .io_d_in_8_a(array_18_io_d_in_8_a),
    .io_d_in_8_valid_a(array_18_io_d_in_8_valid_a),
    .io_d_in_8_b(array_18_io_d_in_8_b),
    .io_d_in_8_valid_b(array_18_io_d_in_8_valid_b),
    .io_d_in_9_a(array_18_io_d_in_9_a),
    .io_d_in_9_valid_a(array_18_io_d_in_9_valid_a),
    .io_d_in_9_b(array_18_io_d_in_9_b),
    .io_d_in_9_valid_b(array_18_io_d_in_9_valid_b),
    .io_d_in_10_a(array_18_io_d_in_10_a),
    .io_d_in_10_valid_a(array_18_io_d_in_10_valid_a),
    .io_d_in_10_b(array_18_io_d_in_10_b),
    .io_d_in_10_valid_b(array_18_io_d_in_10_valid_b),
    .io_d_in_11_a(array_18_io_d_in_11_a),
    .io_d_in_11_valid_a(array_18_io_d_in_11_valid_a),
    .io_d_in_11_b(array_18_io_d_in_11_b),
    .io_d_in_11_valid_b(array_18_io_d_in_11_valid_b),
    .io_d_in_12_a(array_18_io_d_in_12_a),
    .io_d_in_12_valid_a(array_18_io_d_in_12_valid_a),
    .io_d_in_12_b(array_18_io_d_in_12_b),
    .io_d_in_12_valid_b(array_18_io_d_in_12_valid_b),
    .io_d_in_13_a(array_18_io_d_in_13_a),
    .io_d_in_13_valid_a(array_18_io_d_in_13_valid_a),
    .io_d_in_13_b(array_18_io_d_in_13_b),
    .io_d_in_13_valid_b(array_18_io_d_in_13_valid_b),
    .io_d_in_14_a(array_18_io_d_in_14_a),
    .io_d_in_14_valid_a(array_18_io_d_in_14_valid_a),
    .io_d_in_14_b(array_18_io_d_in_14_b),
    .io_d_in_14_valid_b(array_18_io_d_in_14_valid_b),
    .io_d_in_15_a(array_18_io_d_in_15_a),
    .io_d_in_15_valid_a(array_18_io_d_in_15_valid_a),
    .io_d_in_15_b(array_18_io_d_in_15_b),
    .io_d_in_15_valid_b(array_18_io_d_in_15_valid_b),
    .io_d_in_16_a(array_18_io_d_in_16_a),
    .io_d_in_16_valid_a(array_18_io_d_in_16_valid_a),
    .io_d_in_16_b(array_18_io_d_in_16_b),
    .io_d_in_16_valid_b(array_18_io_d_in_16_valid_b),
    .io_d_in_17_a(array_18_io_d_in_17_a),
    .io_d_in_17_valid_a(array_18_io_d_in_17_valid_a),
    .io_d_in_17_b(array_18_io_d_in_17_b),
    .io_d_in_17_valid_b(array_18_io_d_in_17_valid_b),
    .io_d_in_18_a(array_18_io_d_in_18_a),
    .io_d_in_18_valid_a(array_18_io_d_in_18_valid_a),
    .io_d_in_18_b(array_18_io_d_in_18_b),
    .io_d_in_18_valid_b(array_18_io_d_in_18_valid_b),
    .io_d_in_19_a(array_18_io_d_in_19_a),
    .io_d_in_19_valid_a(array_18_io_d_in_19_valid_a),
    .io_d_in_19_b(array_18_io_d_in_19_b),
    .io_d_in_19_valid_b(array_18_io_d_in_19_valid_b),
    .io_d_in_20_a(array_18_io_d_in_20_a),
    .io_d_in_20_valid_a(array_18_io_d_in_20_valid_a),
    .io_d_in_20_b(array_18_io_d_in_20_b),
    .io_d_in_20_valid_b(array_18_io_d_in_20_valid_b),
    .io_d_in_21_a(array_18_io_d_in_21_a),
    .io_d_in_21_valid_a(array_18_io_d_in_21_valid_a),
    .io_d_in_21_b(array_18_io_d_in_21_b),
    .io_d_in_21_valid_b(array_18_io_d_in_21_valid_b),
    .io_d_in_22_a(array_18_io_d_in_22_a),
    .io_d_in_22_valid_a(array_18_io_d_in_22_valid_a),
    .io_d_in_22_b(array_18_io_d_in_22_b),
    .io_d_in_22_valid_b(array_18_io_d_in_22_valid_b),
    .io_d_in_23_a(array_18_io_d_in_23_a),
    .io_d_in_23_valid_a(array_18_io_d_in_23_valid_a),
    .io_d_in_23_b(array_18_io_d_in_23_b),
    .io_d_in_23_valid_b(array_18_io_d_in_23_valid_b),
    .io_d_in_24_a(array_18_io_d_in_24_a),
    .io_d_in_24_valid_a(array_18_io_d_in_24_valid_a),
    .io_d_in_24_b(array_18_io_d_in_24_b),
    .io_d_in_24_valid_b(array_18_io_d_in_24_valid_b),
    .io_d_in_25_a(array_18_io_d_in_25_a),
    .io_d_in_25_valid_a(array_18_io_d_in_25_valid_a),
    .io_d_in_25_b(array_18_io_d_in_25_b),
    .io_d_in_25_valid_b(array_18_io_d_in_25_valid_b),
    .io_d_in_26_a(array_18_io_d_in_26_a),
    .io_d_in_26_valid_a(array_18_io_d_in_26_valid_a),
    .io_d_in_26_b(array_18_io_d_in_26_b),
    .io_d_in_26_valid_b(array_18_io_d_in_26_valid_b),
    .io_d_in_27_a(array_18_io_d_in_27_a),
    .io_d_in_27_valid_a(array_18_io_d_in_27_valid_a),
    .io_d_in_27_b(array_18_io_d_in_27_b),
    .io_d_in_27_valid_b(array_18_io_d_in_27_valid_b),
    .io_d_in_28_a(array_18_io_d_in_28_a),
    .io_d_in_28_valid_a(array_18_io_d_in_28_valid_a),
    .io_d_in_28_b(array_18_io_d_in_28_b),
    .io_d_in_28_valid_b(array_18_io_d_in_28_valid_b),
    .io_d_in_29_a(array_18_io_d_in_29_a),
    .io_d_in_29_valid_a(array_18_io_d_in_29_valid_a),
    .io_d_in_29_b(array_18_io_d_in_29_b),
    .io_d_in_29_valid_b(array_18_io_d_in_29_valid_b),
    .io_d_in_30_a(array_18_io_d_in_30_a),
    .io_d_in_30_valid_a(array_18_io_d_in_30_valid_a),
    .io_d_in_30_b(array_18_io_d_in_30_b),
    .io_d_in_30_valid_b(array_18_io_d_in_30_valid_b),
    .io_d_in_31_a(array_18_io_d_in_31_a),
    .io_d_in_31_valid_a(array_18_io_d_in_31_valid_a),
    .io_d_in_31_b(array_18_io_d_in_31_b),
    .io_d_in_31_valid_b(array_18_io_d_in_31_valid_b),
    .io_d_out_0_a(array_18_io_d_out_0_a),
    .io_d_out_0_valid_a(array_18_io_d_out_0_valid_a),
    .io_d_out_0_b(array_18_io_d_out_0_b),
    .io_d_out_0_valid_b(array_18_io_d_out_0_valid_b),
    .io_d_out_1_a(array_18_io_d_out_1_a),
    .io_d_out_1_valid_a(array_18_io_d_out_1_valid_a),
    .io_d_out_1_b(array_18_io_d_out_1_b),
    .io_d_out_1_valid_b(array_18_io_d_out_1_valid_b),
    .io_d_out_2_a(array_18_io_d_out_2_a),
    .io_d_out_2_valid_a(array_18_io_d_out_2_valid_a),
    .io_d_out_2_b(array_18_io_d_out_2_b),
    .io_d_out_2_valid_b(array_18_io_d_out_2_valid_b),
    .io_d_out_3_a(array_18_io_d_out_3_a),
    .io_d_out_3_valid_a(array_18_io_d_out_3_valid_a),
    .io_d_out_3_b(array_18_io_d_out_3_b),
    .io_d_out_3_valid_b(array_18_io_d_out_3_valid_b),
    .io_d_out_4_a(array_18_io_d_out_4_a),
    .io_d_out_4_valid_a(array_18_io_d_out_4_valid_a),
    .io_d_out_4_b(array_18_io_d_out_4_b),
    .io_d_out_4_valid_b(array_18_io_d_out_4_valid_b),
    .io_d_out_5_a(array_18_io_d_out_5_a),
    .io_d_out_5_valid_a(array_18_io_d_out_5_valid_a),
    .io_d_out_5_b(array_18_io_d_out_5_b),
    .io_d_out_5_valid_b(array_18_io_d_out_5_valid_b),
    .io_d_out_6_a(array_18_io_d_out_6_a),
    .io_d_out_6_valid_a(array_18_io_d_out_6_valid_a),
    .io_d_out_6_b(array_18_io_d_out_6_b),
    .io_d_out_6_valid_b(array_18_io_d_out_6_valid_b),
    .io_d_out_7_a(array_18_io_d_out_7_a),
    .io_d_out_7_valid_a(array_18_io_d_out_7_valid_a),
    .io_d_out_7_b(array_18_io_d_out_7_b),
    .io_d_out_7_valid_b(array_18_io_d_out_7_valid_b),
    .io_d_out_8_a(array_18_io_d_out_8_a),
    .io_d_out_8_valid_a(array_18_io_d_out_8_valid_a),
    .io_d_out_8_b(array_18_io_d_out_8_b),
    .io_d_out_8_valid_b(array_18_io_d_out_8_valid_b),
    .io_d_out_9_a(array_18_io_d_out_9_a),
    .io_d_out_9_valid_a(array_18_io_d_out_9_valid_a),
    .io_d_out_9_b(array_18_io_d_out_9_b),
    .io_d_out_9_valid_b(array_18_io_d_out_9_valid_b),
    .io_d_out_10_a(array_18_io_d_out_10_a),
    .io_d_out_10_valid_a(array_18_io_d_out_10_valid_a),
    .io_d_out_10_b(array_18_io_d_out_10_b),
    .io_d_out_10_valid_b(array_18_io_d_out_10_valid_b),
    .io_d_out_11_a(array_18_io_d_out_11_a),
    .io_d_out_11_valid_a(array_18_io_d_out_11_valid_a),
    .io_d_out_11_b(array_18_io_d_out_11_b),
    .io_d_out_11_valid_b(array_18_io_d_out_11_valid_b),
    .io_d_out_12_a(array_18_io_d_out_12_a),
    .io_d_out_12_valid_a(array_18_io_d_out_12_valid_a),
    .io_d_out_12_b(array_18_io_d_out_12_b),
    .io_d_out_12_valid_b(array_18_io_d_out_12_valid_b),
    .io_d_out_13_a(array_18_io_d_out_13_a),
    .io_d_out_13_valid_a(array_18_io_d_out_13_valid_a),
    .io_d_out_13_b(array_18_io_d_out_13_b),
    .io_d_out_13_valid_b(array_18_io_d_out_13_valid_b),
    .io_d_out_14_a(array_18_io_d_out_14_a),
    .io_d_out_14_valid_a(array_18_io_d_out_14_valid_a),
    .io_d_out_14_b(array_18_io_d_out_14_b),
    .io_d_out_14_valid_b(array_18_io_d_out_14_valid_b),
    .io_d_out_15_a(array_18_io_d_out_15_a),
    .io_d_out_15_valid_a(array_18_io_d_out_15_valid_a),
    .io_d_out_15_b(array_18_io_d_out_15_b),
    .io_d_out_15_valid_b(array_18_io_d_out_15_valid_b),
    .io_d_out_16_a(array_18_io_d_out_16_a),
    .io_d_out_16_valid_a(array_18_io_d_out_16_valid_a),
    .io_d_out_16_b(array_18_io_d_out_16_b),
    .io_d_out_16_valid_b(array_18_io_d_out_16_valid_b),
    .io_d_out_17_a(array_18_io_d_out_17_a),
    .io_d_out_17_valid_a(array_18_io_d_out_17_valid_a),
    .io_d_out_17_b(array_18_io_d_out_17_b),
    .io_d_out_17_valid_b(array_18_io_d_out_17_valid_b),
    .io_d_out_18_a(array_18_io_d_out_18_a),
    .io_d_out_18_valid_a(array_18_io_d_out_18_valid_a),
    .io_d_out_18_b(array_18_io_d_out_18_b),
    .io_d_out_18_valid_b(array_18_io_d_out_18_valid_b),
    .io_d_out_19_a(array_18_io_d_out_19_a),
    .io_d_out_19_valid_a(array_18_io_d_out_19_valid_a),
    .io_d_out_19_b(array_18_io_d_out_19_b),
    .io_d_out_19_valid_b(array_18_io_d_out_19_valid_b),
    .io_d_out_20_a(array_18_io_d_out_20_a),
    .io_d_out_20_valid_a(array_18_io_d_out_20_valid_a),
    .io_d_out_20_b(array_18_io_d_out_20_b),
    .io_d_out_20_valid_b(array_18_io_d_out_20_valid_b),
    .io_d_out_21_a(array_18_io_d_out_21_a),
    .io_d_out_21_valid_a(array_18_io_d_out_21_valid_a),
    .io_d_out_21_b(array_18_io_d_out_21_b),
    .io_d_out_21_valid_b(array_18_io_d_out_21_valid_b),
    .io_d_out_22_a(array_18_io_d_out_22_a),
    .io_d_out_22_valid_a(array_18_io_d_out_22_valid_a),
    .io_d_out_22_b(array_18_io_d_out_22_b),
    .io_d_out_22_valid_b(array_18_io_d_out_22_valid_b),
    .io_d_out_23_a(array_18_io_d_out_23_a),
    .io_d_out_23_valid_a(array_18_io_d_out_23_valid_a),
    .io_d_out_23_b(array_18_io_d_out_23_b),
    .io_d_out_23_valid_b(array_18_io_d_out_23_valid_b),
    .io_d_out_24_a(array_18_io_d_out_24_a),
    .io_d_out_24_valid_a(array_18_io_d_out_24_valid_a),
    .io_d_out_24_b(array_18_io_d_out_24_b),
    .io_d_out_24_valid_b(array_18_io_d_out_24_valid_b),
    .io_d_out_25_a(array_18_io_d_out_25_a),
    .io_d_out_25_valid_a(array_18_io_d_out_25_valid_a),
    .io_d_out_25_b(array_18_io_d_out_25_b),
    .io_d_out_25_valid_b(array_18_io_d_out_25_valid_b),
    .io_d_out_26_a(array_18_io_d_out_26_a),
    .io_d_out_26_valid_a(array_18_io_d_out_26_valid_a),
    .io_d_out_26_b(array_18_io_d_out_26_b),
    .io_d_out_26_valid_b(array_18_io_d_out_26_valid_b),
    .io_d_out_27_a(array_18_io_d_out_27_a),
    .io_d_out_27_valid_a(array_18_io_d_out_27_valid_a),
    .io_d_out_27_b(array_18_io_d_out_27_b),
    .io_d_out_27_valid_b(array_18_io_d_out_27_valid_b),
    .io_d_out_28_a(array_18_io_d_out_28_a),
    .io_d_out_28_valid_a(array_18_io_d_out_28_valid_a),
    .io_d_out_28_b(array_18_io_d_out_28_b),
    .io_d_out_28_valid_b(array_18_io_d_out_28_valid_b),
    .io_d_out_29_a(array_18_io_d_out_29_a),
    .io_d_out_29_valid_a(array_18_io_d_out_29_valid_a),
    .io_d_out_29_b(array_18_io_d_out_29_b),
    .io_d_out_29_valid_b(array_18_io_d_out_29_valid_b),
    .io_d_out_30_a(array_18_io_d_out_30_a),
    .io_d_out_30_valid_a(array_18_io_d_out_30_valid_a),
    .io_d_out_30_b(array_18_io_d_out_30_b),
    .io_d_out_30_valid_b(array_18_io_d_out_30_valid_b),
    .io_d_out_31_a(array_18_io_d_out_31_a),
    .io_d_out_31_valid_a(array_18_io_d_out_31_valid_a),
    .io_d_out_31_b(array_18_io_d_out_31_b),
    .io_d_out_31_valid_b(array_18_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_18_io_wr_en_mem1),
    .io_wr_en_mem2(array_18_io_wr_en_mem2),
    .io_wr_en_mem3(array_18_io_wr_en_mem3),
    .io_wr_en_mem4(array_18_io_wr_en_mem4),
    .io_wr_en_mem5(array_18_io_wr_en_mem5),
    .io_wr_en_mem6(array_18_io_wr_en_mem6),
    .io_wr_instr_mem1(array_18_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_18_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_18_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_18_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_18_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_18_io_wr_instr_mem6),
    .io_PC1_in(array_18_io_PC1_in),
    .io_PC6_out(array_18_io_PC6_out),
    .io_Addr_in(array_18_io_Addr_in),
    .io_Addr_out(array_18_io_Addr_out)
  );
  BuildingBlockNew array_19 ( // @[BP.scala 45:51]
    .clock(array_19_clock),
    .reset(array_19_reset),
    .io_d_in_0_a(array_19_io_d_in_0_a),
    .io_d_in_0_valid_a(array_19_io_d_in_0_valid_a),
    .io_d_in_0_b(array_19_io_d_in_0_b),
    .io_d_in_0_valid_b(array_19_io_d_in_0_valid_b),
    .io_d_in_1_a(array_19_io_d_in_1_a),
    .io_d_in_1_valid_a(array_19_io_d_in_1_valid_a),
    .io_d_in_1_b(array_19_io_d_in_1_b),
    .io_d_in_1_valid_b(array_19_io_d_in_1_valid_b),
    .io_d_in_2_a(array_19_io_d_in_2_a),
    .io_d_in_2_valid_a(array_19_io_d_in_2_valid_a),
    .io_d_in_2_b(array_19_io_d_in_2_b),
    .io_d_in_2_valid_b(array_19_io_d_in_2_valid_b),
    .io_d_in_3_a(array_19_io_d_in_3_a),
    .io_d_in_3_valid_a(array_19_io_d_in_3_valid_a),
    .io_d_in_3_b(array_19_io_d_in_3_b),
    .io_d_in_3_valid_b(array_19_io_d_in_3_valid_b),
    .io_d_in_4_a(array_19_io_d_in_4_a),
    .io_d_in_4_valid_a(array_19_io_d_in_4_valid_a),
    .io_d_in_4_b(array_19_io_d_in_4_b),
    .io_d_in_4_valid_b(array_19_io_d_in_4_valid_b),
    .io_d_in_5_a(array_19_io_d_in_5_a),
    .io_d_in_5_valid_a(array_19_io_d_in_5_valid_a),
    .io_d_in_5_b(array_19_io_d_in_5_b),
    .io_d_in_5_valid_b(array_19_io_d_in_5_valid_b),
    .io_d_in_6_a(array_19_io_d_in_6_a),
    .io_d_in_6_valid_a(array_19_io_d_in_6_valid_a),
    .io_d_in_6_b(array_19_io_d_in_6_b),
    .io_d_in_6_valid_b(array_19_io_d_in_6_valid_b),
    .io_d_in_7_a(array_19_io_d_in_7_a),
    .io_d_in_7_valid_a(array_19_io_d_in_7_valid_a),
    .io_d_in_7_b(array_19_io_d_in_7_b),
    .io_d_in_7_valid_b(array_19_io_d_in_7_valid_b),
    .io_d_in_8_a(array_19_io_d_in_8_a),
    .io_d_in_8_valid_a(array_19_io_d_in_8_valid_a),
    .io_d_in_8_b(array_19_io_d_in_8_b),
    .io_d_in_8_valid_b(array_19_io_d_in_8_valid_b),
    .io_d_in_9_a(array_19_io_d_in_9_a),
    .io_d_in_9_valid_a(array_19_io_d_in_9_valid_a),
    .io_d_in_9_b(array_19_io_d_in_9_b),
    .io_d_in_9_valid_b(array_19_io_d_in_9_valid_b),
    .io_d_in_10_a(array_19_io_d_in_10_a),
    .io_d_in_10_valid_a(array_19_io_d_in_10_valid_a),
    .io_d_in_10_b(array_19_io_d_in_10_b),
    .io_d_in_10_valid_b(array_19_io_d_in_10_valid_b),
    .io_d_in_11_a(array_19_io_d_in_11_a),
    .io_d_in_11_valid_a(array_19_io_d_in_11_valid_a),
    .io_d_in_11_b(array_19_io_d_in_11_b),
    .io_d_in_11_valid_b(array_19_io_d_in_11_valid_b),
    .io_d_in_12_a(array_19_io_d_in_12_a),
    .io_d_in_12_valid_a(array_19_io_d_in_12_valid_a),
    .io_d_in_12_b(array_19_io_d_in_12_b),
    .io_d_in_12_valid_b(array_19_io_d_in_12_valid_b),
    .io_d_in_13_a(array_19_io_d_in_13_a),
    .io_d_in_13_valid_a(array_19_io_d_in_13_valid_a),
    .io_d_in_13_b(array_19_io_d_in_13_b),
    .io_d_in_13_valid_b(array_19_io_d_in_13_valid_b),
    .io_d_in_14_a(array_19_io_d_in_14_a),
    .io_d_in_14_valid_a(array_19_io_d_in_14_valid_a),
    .io_d_in_14_b(array_19_io_d_in_14_b),
    .io_d_in_14_valid_b(array_19_io_d_in_14_valid_b),
    .io_d_in_15_a(array_19_io_d_in_15_a),
    .io_d_in_15_valid_a(array_19_io_d_in_15_valid_a),
    .io_d_in_15_b(array_19_io_d_in_15_b),
    .io_d_in_15_valid_b(array_19_io_d_in_15_valid_b),
    .io_d_in_16_a(array_19_io_d_in_16_a),
    .io_d_in_16_valid_a(array_19_io_d_in_16_valid_a),
    .io_d_in_16_b(array_19_io_d_in_16_b),
    .io_d_in_16_valid_b(array_19_io_d_in_16_valid_b),
    .io_d_in_17_a(array_19_io_d_in_17_a),
    .io_d_in_17_valid_a(array_19_io_d_in_17_valid_a),
    .io_d_in_17_b(array_19_io_d_in_17_b),
    .io_d_in_17_valid_b(array_19_io_d_in_17_valid_b),
    .io_d_in_18_a(array_19_io_d_in_18_a),
    .io_d_in_18_valid_a(array_19_io_d_in_18_valid_a),
    .io_d_in_18_b(array_19_io_d_in_18_b),
    .io_d_in_18_valid_b(array_19_io_d_in_18_valid_b),
    .io_d_in_19_a(array_19_io_d_in_19_a),
    .io_d_in_19_valid_a(array_19_io_d_in_19_valid_a),
    .io_d_in_19_b(array_19_io_d_in_19_b),
    .io_d_in_19_valid_b(array_19_io_d_in_19_valid_b),
    .io_d_in_20_a(array_19_io_d_in_20_a),
    .io_d_in_20_valid_a(array_19_io_d_in_20_valid_a),
    .io_d_in_20_b(array_19_io_d_in_20_b),
    .io_d_in_20_valid_b(array_19_io_d_in_20_valid_b),
    .io_d_in_21_a(array_19_io_d_in_21_a),
    .io_d_in_21_valid_a(array_19_io_d_in_21_valid_a),
    .io_d_in_21_b(array_19_io_d_in_21_b),
    .io_d_in_21_valid_b(array_19_io_d_in_21_valid_b),
    .io_d_in_22_a(array_19_io_d_in_22_a),
    .io_d_in_22_valid_a(array_19_io_d_in_22_valid_a),
    .io_d_in_22_b(array_19_io_d_in_22_b),
    .io_d_in_22_valid_b(array_19_io_d_in_22_valid_b),
    .io_d_in_23_a(array_19_io_d_in_23_a),
    .io_d_in_23_valid_a(array_19_io_d_in_23_valid_a),
    .io_d_in_23_b(array_19_io_d_in_23_b),
    .io_d_in_23_valid_b(array_19_io_d_in_23_valid_b),
    .io_d_in_24_a(array_19_io_d_in_24_a),
    .io_d_in_24_valid_a(array_19_io_d_in_24_valid_a),
    .io_d_in_24_b(array_19_io_d_in_24_b),
    .io_d_in_24_valid_b(array_19_io_d_in_24_valid_b),
    .io_d_in_25_a(array_19_io_d_in_25_a),
    .io_d_in_25_valid_a(array_19_io_d_in_25_valid_a),
    .io_d_in_25_b(array_19_io_d_in_25_b),
    .io_d_in_25_valid_b(array_19_io_d_in_25_valid_b),
    .io_d_in_26_a(array_19_io_d_in_26_a),
    .io_d_in_26_valid_a(array_19_io_d_in_26_valid_a),
    .io_d_in_26_b(array_19_io_d_in_26_b),
    .io_d_in_26_valid_b(array_19_io_d_in_26_valid_b),
    .io_d_in_27_a(array_19_io_d_in_27_a),
    .io_d_in_27_valid_a(array_19_io_d_in_27_valid_a),
    .io_d_in_27_b(array_19_io_d_in_27_b),
    .io_d_in_27_valid_b(array_19_io_d_in_27_valid_b),
    .io_d_in_28_a(array_19_io_d_in_28_a),
    .io_d_in_28_valid_a(array_19_io_d_in_28_valid_a),
    .io_d_in_28_b(array_19_io_d_in_28_b),
    .io_d_in_28_valid_b(array_19_io_d_in_28_valid_b),
    .io_d_in_29_a(array_19_io_d_in_29_a),
    .io_d_in_29_valid_a(array_19_io_d_in_29_valid_a),
    .io_d_in_29_b(array_19_io_d_in_29_b),
    .io_d_in_29_valid_b(array_19_io_d_in_29_valid_b),
    .io_d_in_30_a(array_19_io_d_in_30_a),
    .io_d_in_30_valid_a(array_19_io_d_in_30_valid_a),
    .io_d_in_30_b(array_19_io_d_in_30_b),
    .io_d_in_30_valid_b(array_19_io_d_in_30_valid_b),
    .io_d_in_31_a(array_19_io_d_in_31_a),
    .io_d_in_31_valid_a(array_19_io_d_in_31_valid_a),
    .io_d_in_31_b(array_19_io_d_in_31_b),
    .io_d_in_31_valid_b(array_19_io_d_in_31_valid_b),
    .io_d_out_0_a(array_19_io_d_out_0_a),
    .io_d_out_0_valid_a(array_19_io_d_out_0_valid_a),
    .io_d_out_0_b(array_19_io_d_out_0_b),
    .io_d_out_0_valid_b(array_19_io_d_out_0_valid_b),
    .io_d_out_1_a(array_19_io_d_out_1_a),
    .io_d_out_1_valid_a(array_19_io_d_out_1_valid_a),
    .io_d_out_1_b(array_19_io_d_out_1_b),
    .io_d_out_1_valid_b(array_19_io_d_out_1_valid_b),
    .io_d_out_2_a(array_19_io_d_out_2_a),
    .io_d_out_2_valid_a(array_19_io_d_out_2_valid_a),
    .io_d_out_2_b(array_19_io_d_out_2_b),
    .io_d_out_2_valid_b(array_19_io_d_out_2_valid_b),
    .io_d_out_3_a(array_19_io_d_out_3_a),
    .io_d_out_3_valid_a(array_19_io_d_out_3_valid_a),
    .io_d_out_3_b(array_19_io_d_out_3_b),
    .io_d_out_3_valid_b(array_19_io_d_out_3_valid_b),
    .io_d_out_4_a(array_19_io_d_out_4_a),
    .io_d_out_4_valid_a(array_19_io_d_out_4_valid_a),
    .io_d_out_4_b(array_19_io_d_out_4_b),
    .io_d_out_4_valid_b(array_19_io_d_out_4_valid_b),
    .io_d_out_5_a(array_19_io_d_out_5_a),
    .io_d_out_5_valid_a(array_19_io_d_out_5_valid_a),
    .io_d_out_5_b(array_19_io_d_out_5_b),
    .io_d_out_5_valid_b(array_19_io_d_out_5_valid_b),
    .io_d_out_6_a(array_19_io_d_out_6_a),
    .io_d_out_6_valid_a(array_19_io_d_out_6_valid_a),
    .io_d_out_6_b(array_19_io_d_out_6_b),
    .io_d_out_6_valid_b(array_19_io_d_out_6_valid_b),
    .io_d_out_7_a(array_19_io_d_out_7_a),
    .io_d_out_7_valid_a(array_19_io_d_out_7_valid_a),
    .io_d_out_7_b(array_19_io_d_out_7_b),
    .io_d_out_7_valid_b(array_19_io_d_out_7_valid_b),
    .io_d_out_8_a(array_19_io_d_out_8_a),
    .io_d_out_8_valid_a(array_19_io_d_out_8_valid_a),
    .io_d_out_8_b(array_19_io_d_out_8_b),
    .io_d_out_8_valid_b(array_19_io_d_out_8_valid_b),
    .io_d_out_9_a(array_19_io_d_out_9_a),
    .io_d_out_9_valid_a(array_19_io_d_out_9_valid_a),
    .io_d_out_9_b(array_19_io_d_out_9_b),
    .io_d_out_9_valid_b(array_19_io_d_out_9_valid_b),
    .io_d_out_10_a(array_19_io_d_out_10_a),
    .io_d_out_10_valid_a(array_19_io_d_out_10_valid_a),
    .io_d_out_10_b(array_19_io_d_out_10_b),
    .io_d_out_10_valid_b(array_19_io_d_out_10_valid_b),
    .io_d_out_11_a(array_19_io_d_out_11_a),
    .io_d_out_11_valid_a(array_19_io_d_out_11_valid_a),
    .io_d_out_11_b(array_19_io_d_out_11_b),
    .io_d_out_11_valid_b(array_19_io_d_out_11_valid_b),
    .io_d_out_12_a(array_19_io_d_out_12_a),
    .io_d_out_12_valid_a(array_19_io_d_out_12_valid_a),
    .io_d_out_12_b(array_19_io_d_out_12_b),
    .io_d_out_12_valid_b(array_19_io_d_out_12_valid_b),
    .io_d_out_13_a(array_19_io_d_out_13_a),
    .io_d_out_13_valid_a(array_19_io_d_out_13_valid_a),
    .io_d_out_13_b(array_19_io_d_out_13_b),
    .io_d_out_13_valid_b(array_19_io_d_out_13_valid_b),
    .io_d_out_14_a(array_19_io_d_out_14_a),
    .io_d_out_14_valid_a(array_19_io_d_out_14_valid_a),
    .io_d_out_14_b(array_19_io_d_out_14_b),
    .io_d_out_14_valid_b(array_19_io_d_out_14_valid_b),
    .io_d_out_15_a(array_19_io_d_out_15_a),
    .io_d_out_15_valid_a(array_19_io_d_out_15_valid_a),
    .io_d_out_15_b(array_19_io_d_out_15_b),
    .io_d_out_15_valid_b(array_19_io_d_out_15_valid_b),
    .io_d_out_16_a(array_19_io_d_out_16_a),
    .io_d_out_16_valid_a(array_19_io_d_out_16_valid_a),
    .io_d_out_16_b(array_19_io_d_out_16_b),
    .io_d_out_16_valid_b(array_19_io_d_out_16_valid_b),
    .io_d_out_17_a(array_19_io_d_out_17_a),
    .io_d_out_17_valid_a(array_19_io_d_out_17_valid_a),
    .io_d_out_17_b(array_19_io_d_out_17_b),
    .io_d_out_17_valid_b(array_19_io_d_out_17_valid_b),
    .io_d_out_18_a(array_19_io_d_out_18_a),
    .io_d_out_18_valid_a(array_19_io_d_out_18_valid_a),
    .io_d_out_18_b(array_19_io_d_out_18_b),
    .io_d_out_18_valid_b(array_19_io_d_out_18_valid_b),
    .io_d_out_19_a(array_19_io_d_out_19_a),
    .io_d_out_19_valid_a(array_19_io_d_out_19_valid_a),
    .io_d_out_19_b(array_19_io_d_out_19_b),
    .io_d_out_19_valid_b(array_19_io_d_out_19_valid_b),
    .io_d_out_20_a(array_19_io_d_out_20_a),
    .io_d_out_20_valid_a(array_19_io_d_out_20_valid_a),
    .io_d_out_20_b(array_19_io_d_out_20_b),
    .io_d_out_20_valid_b(array_19_io_d_out_20_valid_b),
    .io_d_out_21_a(array_19_io_d_out_21_a),
    .io_d_out_21_valid_a(array_19_io_d_out_21_valid_a),
    .io_d_out_21_b(array_19_io_d_out_21_b),
    .io_d_out_21_valid_b(array_19_io_d_out_21_valid_b),
    .io_d_out_22_a(array_19_io_d_out_22_a),
    .io_d_out_22_valid_a(array_19_io_d_out_22_valid_a),
    .io_d_out_22_b(array_19_io_d_out_22_b),
    .io_d_out_22_valid_b(array_19_io_d_out_22_valid_b),
    .io_d_out_23_a(array_19_io_d_out_23_a),
    .io_d_out_23_valid_a(array_19_io_d_out_23_valid_a),
    .io_d_out_23_b(array_19_io_d_out_23_b),
    .io_d_out_23_valid_b(array_19_io_d_out_23_valid_b),
    .io_d_out_24_a(array_19_io_d_out_24_a),
    .io_d_out_24_valid_a(array_19_io_d_out_24_valid_a),
    .io_d_out_24_b(array_19_io_d_out_24_b),
    .io_d_out_24_valid_b(array_19_io_d_out_24_valid_b),
    .io_d_out_25_a(array_19_io_d_out_25_a),
    .io_d_out_25_valid_a(array_19_io_d_out_25_valid_a),
    .io_d_out_25_b(array_19_io_d_out_25_b),
    .io_d_out_25_valid_b(array_19_io_d_out_25_valid_b),
    .io_d_out_26_a(array_19_io_d_out_26_a),
    .io_d_out_26_valid_a(array_19_io_d_out_26_valid_a),
    .io_d_out_26_b(array_19_io_d_out_26_b),
    .io_d_out_26_valid_b(array_19_io_d_out_26_valid_b),
    .io_d_out_27_a(array_19_io_d_out_27_a),
    .io_d_out_27_valid_a(array_19_io_d_out_27_valid_a),
    .io_d_out_27_b(array_19_io_d_out_27_b),
    .io_d_out_27_valid_b(array_19_io_d_out_27_valid_b),
    .io_d_out_28_a(array_19_io_d_out_28_a),
    .io_d_out_28_valid_a(array_19_io_d_out_28_valid_a),
    .io_d_out_28_b(array_19_io_d_out_28_b),
    .io_d_out_28_valid_b(array_19_io_d_out_28_valid_b),
    .io_d_out_29_a(array_19_io_d_out_29_a),
    .io_d_out_29_valid_a(array_19_io_d_out_29_valid_a),
    .io_d_out_29_b(array_19_io_d_out_29_b),
    .io_d_out_29_valid_b(array_19_io_d_out_29_valid_b),
    .io_d_out_30_a(array_19_io_d_out_30_a),
    .io_d_out_30_valid_a(array_19_io_d_out_30_valid_a),
    .io_d_out_30_b(array_19_io_d_out_30_b),
    .io_d_out_30_valid_b(array_19_io_d_out_30_valid_b),
    .io_d_out_31_a(array_19_io_d_out_31_a),
    .io_d_out_31_valid_a(array_19_io_d_out_31_valid_a),
    .io_d_out_31_b(array_19_io_d_out_31_b),
    .io_d_out_31_valid_b(array_19_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_19_io_wr_en_mem1),
    .io_wr_en_mem2(array_19_io_wr_en_mem2),
    .io_wr_en_mem3(array_19_io_wr_en_mem3),
    .io_wr_en_mem4(array_19_io_wr_en_mem4),
    .io_wr_en_mem5(array_19_io_wr_en_mem5),
    .io_wr_en_mem6(array_19_io_wr_en_mem6),
    .io_wr_instr_mem1(array_19_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_19_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_19_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_19_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_19_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_19_io_wr_instr_mem6),
    .io_PC1_in(array_19_io_PC1_in),
    .io_PC6_out(array_19_io_PC6_out),
    .io_Addr_in(array_19_io_Addr_in),
    .io_Addr_out(array_19_io_Addr_out)
  );
  BuildingBlockNew array_20 ( // @[BP.scala 45:51]
    .clock(array_20_clock),
    .reset(array_20_reset),
    .io_d_in_0_a(array_20_io_d_in_0_a),
    .io_d_in_0_valid_a(array_20_io_d_in_0_valid_a),
    .io_d_in_0_b(array_20_io_d_in_0_b),
    .io_d_in_0_valid_b(array_20_io_d_in_0_valid_b),
    .io_d_in_1_a(array_20_io_d_in_1_a),
    .io_d_in_1_valid_a(array_20_io_d_in_1_valid_a),
    .io_d_in_1_b(array_20_io_d_in_1_b),
    .io_d_in_1_valid_b(array_20_io_d_in_1_valid_b),
    .io_d_in_2_a(array_20_io_d_in_2_a),
    .io_d_in_2_valid_a(array_20_io_d_in_2_valid_a),
    .io_d_in_2_b(array_20_io_d_in_2_b),
    .io_d_in_2_valid_b(array_20_io_d_in_2_valid_b),
    .io_d_in_3_a(array_20_io_d_in_3_a),
    .io_d_in_3_valid_a(array_20_io_d_in_3_valid_a),
    .io_d_in_3_b(array_20_io_d_in_3_b),
    .io_d_in_3_valid_b(array_20_io_d_in_3_valid_b),
    .io_d_in_4_a(array_20_io_d_in_4_a),
    .io_d_in_4_valid_a(array_20_io_d_in_4_valid_a),
    .io_d_in_4_b(array_20_io_d_in_4_b),
    .io_d_in_4_valid_b(array_20_io_d_in_4_valid_b),
    .io_d_in_5_a(array_20_io_d_in_5_a),
    .io_d_in_5_valid_a(array_20_io_d_in_5_valid_a),
    .io_d_in_5_b(array_20_io_d_in_5_b),
    .io_d_in_5_valid_b(array_20_io_d_in_5_valid_b),
    .io_d_in_6_a(array_20_io_d_in_6_a),
    .io_d_in_6_valid_a(array_20_io_d_in_6_valid_a),
    .io_d_in_6_b(array_20_io_d_in_6_b),
    .io_d_in_6_valid_b(array_20_io_d_in_6_valid_b),
    .io_d_in_7_a(array_20_io_d_in_7_a),
    .io_d_in_7_valid_a(array_20_io_d_in_7_valid_a),
    .io_d_in_7_b(array_20_io_d_in_7_b),
    .io_d_in_7_valid_b(array_20_io_d_in_7_valid_b),
    .io_d_in_8_a(array_20_io_d_in_8_a),
    .io_d_in_8_valid_a(array_20_io_d_in_8_valid_a),
    .io_d_in_8_b(array_20_io_d_in_8_b),
    .io_d_in_8_valid_b(array_20_io_d_in_8_valid_b),
    .io_d_in_9_a(array_20_io_d_in_9_a),
    .io_d_in_9_valid_a(array_20_io_d_in_9_valid_a),
    .io_d_in_9_b(array_20_io_d_in_9_b),
    .io_d_in_9_valid_b(array_20_io_d_in_9_valid_b),
    .io_d_in_10_a(array_20_io_d_in_10_a),
    .io_d_in_10_valid_a(array_20_io_d_in_10_valid_a),
    .io_d_in_10_b(array_20_io_d_in_10_b),
    .io_d_in_10_valid_b(array_20_io_d_in_10_valid_b),
    .io_d_in_11_a(array_20_io_d_in_11_a),
    .io_d_in_11_valid_a(array_20_io_d_in_11_valid_a),
    .io_d_in_11_b(array_20_io_d_in_11_b),
    .io_d_in_11_valid_b(array_20_io_d_in_11_valid_b),
    .io_d_in_12_a(array_20_io_d_in_12_a),
    .io_d_in_12_valid_a(array_20_io_d_in_12_valid_a),
    .io_d_in_12_b(array_20_io_d_in_12_b),
    .io_d_in_12_valid_b(array_20_io_d_in_12_valid_b),
    .io_d_in_13_a(array_20_io_d_in_13_a),
    .io_d_in_13_valid_a(array_20_io_d_in_13_valid_a),
    .io_d_in_13_b(array_20_io_d_in_13_b),
    .io_d_in_13_valid_b(array_20_io_d_in_13_valid_b),
    .io_d_in_14_a(array_20_io_d_in_14_a),
    .io_d_in_14_valid_a(array_20_io_d_in_14_valid_a),
    .io_d_in_14_b(array_20_io_d_in_14_b),
    .io_d_in_14_valid_b(array_20_io_d_in_14_valid_b),
    .io_d_in_15_a(array_20_io_d_in_15_a),
    .io_d_in_15_valid_a(array_20_io_d_in_15_valid_a),
    .io_d_in_15_b(array_20_io_d_in_15_b),
    .io_d_in_15_valid_b(array_20_io_d_in_15_valid_b),
    .io_d_in_16_a(array_20_io_d_in_16_a),
    .io_d_in_16_valid_a(array_20_io_d_in_16_valid_a),
    .io_d_in_16_b(array_20_io_d_in_16_b),
    .io_d_in_16_valid_b(array_20_io_d_in_16_valid_b),
    .io_d_in_17_a(array_20_io_d_in_17_a),
    .io_d_in_17_valid_a(array_20_io_d_in_17_valid_a),
    .io_d_in_17_b(array_20_io_d_in_17_b),
    .io_d_in_17_valid_b(array_20_io_d_in_17_valid_b),
    .io_d_in_18_a(array_20_io_d_in_18_a),
    .io_d_in_18_valid_a(array_20_io_d_in_18_valid_a),
    .io_d_in_18_b(array_20_io_d_in_18_b),
    .io_d_in_18_valid_b(array_20_io_d_in_18_valid_b),
    .io_d_in_19_a(array_20_io_d_in_19_a),
    .io_d_in_19_valid_a(array_20_io_d_in_19_valid_a),
    .io_d_in_19_b(array_20_io_d_in_19_b),
    .io_d_in_19_valid_b(array_20_io_d_in_19_valid_b),
    .io_d_in_20_a(array_20_io_d_in_20_a),
    .io_d_in_20_valid_a(array_20_io_d_in_20_valid_a),
    .io_d_in_20_b(array_20_io_d_in_20_b),
    .io_d_in_20_valid_b(array_20_io_d_in_20_valid_b),
    .io_d_in_21_a(array_20_io_d_in_21_a),
    .io_d_in_21_valid_a(array_20_io_d_in_21_valid_a),
    .io_d_in_21_b(array_20_io_d_in_21_b),
    .io_d_in_21_valid_b(array_20_io_d_in_21_valid_b),
    .io_d_in_22_a(array_20_io_d_in_22_a),
    .io_d_in_22_valid_a(array_20_io_d_in_22_valid_a),
    .io_d_in_22_b(array_20_io_d_in_22_b),
    .io_d_in_22_valid_b(array_20_io_d_in_22_valid_b),
    .io_d_in_23_a(array_20_io_d_in_23_a),
    .io_d_in_23_valid_a(array_20_io_d_in_23_valid_a),
    .io_d_in_23_b(array_20_io_d_in_23_b),
    .io_d_in_23_valid_b(array_20_io_d_in_23_valid_b),
    .io_d_in_24_a(array_20_io_d_in_24_a),
    .io_d_in_24_valid_a(array_20_io_d_in_24_valid_a),
    .io_d_in_24_b(array_20_io_d_in_24_b),
    .io_d_in_24_valid_b(array_20_io_d_in_24_valid_b),
    .io_d_in_25_a(array_20_io_d_in_25_a),
    .io_d_in_25_valid_a(array_20_io_d_in_25_valid_a),
    .io_d_in_25_b(array_20_io_d_in_25_b),
    .io_d_in_25_valid_b(array_20_io_d_in_25_valid_b),
    .io_d_in_26_a(array_20_io_d_in_26_a),
    .io_d_in_26_valid_a(array_20_io_d_in_26_valid_a),
    .io_d_in_26_b(array_20_io_d_in_26_b),
    .io_d_in_26_valid_b(array_20_io_d_in_26_valid_b),
    .io_d_in_27_a(array_20_io_d_in_27_a),
    .io_d_in_27_valid_a(array_20_io_d_in_27_valid_a),
    .io_d_in_27_b(array_20_io_d_in_27_b),
    .io_d_in_27_valid_b(array_20_io_d_in_27_valid_b),
    .io_d_in_28_a(array_20_io_d_in_28_a),
    .io_d_in_28_valid_a(array_20_io_d_in_28_valid_a),
    .io_d_in_28_b(array_20_io_d_in_28_b),
    .io_d_in_28_valid_b(array_20_io_d_in_28_valid_b),
    .io_d_in_29_a(array_20_io_d_in_29_a),
    .io_d_in_29_valid_a(array_20_io_d_in_29_valid_a),
    .io_d_in_29_b(array_20_io_d_in_29_b),
    .io_d_in_29_valid_b(array_20_io_d_in_29_valid_b),
    .io_d_in_30_a(array_20_io_d_in_30_a),
    .io_d_in_30_valid_a(array_20_io_d_in_30_valid_a),
    .io_d_in_30_b(array_20_io_d_in_30_b),
    .io_d_in_30_valid_b(array_20_io_d_in_30_valid_b),
    .io_d_in_31_a(array_20_io_d_in_31_a),
    .io_d_in_31_valid_a(array_20_io_d_in_31_valid_a),
    .io_d_in_31_b(array_20_io_d_in_31_b),
    .io_d_in_31_valid_b(array_20_io_d_in_31_valid_b),
    .io_d_out_0_a(array_20_io_d_out_0_a),
    .io_d_out_0_valid_a(array_20_io_d_out_0_valid_a),
    .io_d_out_0_b(array_20_io_d_out_0_b),
    .io_d_out_0_valid_b(array_20_io_d_out_0_valid_b),
    .io_d_out_1_a(array_20_io_d_out_1_a),
    .io_d_out_1_valid_a(array_20_io_d_out_1_valid_a),
    .io_d_out_1_b(array_20_io_d_out_1_b),
    .io_d_out_1_valid_b(array_20_io_d_out_1_valid_b),
    .io_d_out_2_a(array_20_io_d_out_2_a),
    .io_d_out_2_valid_a(array_20_io_d_out_2_valid_a),
    .io_d_out_2_b(array_20_io_d_out_2_b),
    .io_d_out_2_valid_b(array_20_io_d_out_2_valid_b),
    .io_d_out_3_a(array_20_io_d_out_3_a),
    .io_d_out_3_valid_a(array_20_io_d_out_3_valid_a),
    .io_d_out_3_b(array_20_io_d_out_3_b),
    .io_d_out_3_valid_b(array_20_io_d_out_3_valid_b),
    .io_d_out_4_a(array_20_io_d_out_4_a),
    .io_d_out_4_valid_a(array_20_io_d_out_4_valid_a),
    .io_d_out_4_b(array_20_io_d_out_4_b),
    .io_d_out_4_valid_b(array_20_io_d_out_4_valid_b),
    .io_d_out_5_a(array_20_io_d_out_5_a),
    .io_d_out_5_valid_a(array_20_io_d_out_5_valid_a),
    .io_d_out_5_b(array_20_io_d_out_5_b),
    .io_d_out_5_valid_b(array_20_io_d_out_5_valid_b),
    .io_d_out_6_a(array_20_io_d_out_6_a),
    .io_d_out_6_valid_a(array_20_io_d_out_6_valid_a),
    .io_d_out_6_b(array_20_io_d_out_6_b),
    .io_d_out_6_valid_b(array_20_io_d_out_6_valid_b),
    .io_d_out_7_a(array_20_io_d_out_7_a),
    .io_d_out_7_valid_a(array_20_io_d_out_7_valid_a),
    .io_d_out_7_b(array_20_io_d_out_7_b),
    .io_d_out_7_valid_b(array_20_io_d_out_7_valid_b),
    .io_d_out_8_a(array_20_io_d_out_8_a),
    .io_d_out_8_valid_a(array_20_io_d_out_8_valid_a),
    .io_d_out_8_b(array_20_io_d_out_8_b),
    .io_d_out_8_valid_b(array_20_io_d_out_8_valid_b),
    .io_d_out_9_a(array_20_io_d_out_9_a),
    .io_d_out_9_valid_a(array_20_io_d_out_9_valid_a),
    .io_d_out_9_b(array_20_io_d_out_9_b),
    .io_d_out_9_valid_b(array_20_io_d_out_9_valid_b),
    .io_d_out_10_a(array_20_io_d_out_10_a),
    .io_d_out_10_valid_a(array_20_io_d_out_10_valid_a),
    .io_d_out_10_b(array_20_io_d_out_10_b),
    .io_d_out_10_valid_b(array_20_io_d_out_10_valid_b),
    .io_d_out_11_a(array_20_io_d_out_11_a),
    .io_d_out_11_valid_a(array_20_io_d_out_11_valid_a),
    .io_d_out_11_b(array_20_io_d_out_11_b),
    .io_d_out_11_valid_b(array_20_io_d_out_11_valid_b),
    .io_d_out_12_a(array_20_io_d_out_12_a),
    .io_d_out_12_valid_a(array_20_io_d_out_12_valid_a),
    .io_d_out_12_b(array_20_io_d_out_12_b),
    .io_d_out_12_valid_b(array_20_io_d_out_12_valid_b),
    .io_d_out_13_a(array_20_io_d_out_13_a),
    .io_d_out_13_valid_a(array_20_io_d_out_13_valid_a),
    .io_d_out_13_b(array_20_io_d_out_13_b),
    .io_d_out_13_valid_b(array_20_io_d_out_13_valid_b),
    .io_d_out_14_a(array_20_io_d_out_14_a),
    .io_d_out_14_valid_a(array_20_io_d_out_14_valid_a),
    .io_d_out_14_b(array_20_io_d_out_14_b),
    .io_d_out_14_valid_b(array_20_io_d_out_14_valid_b),
    .io_d_out_15_a(array_20_io_d_out_15_a),
    .io_d_out_15_valid_a(array_20_io_d_out_15_valid_a),
    .io_d_out_15_b(array_20_io_d_out_15_b),
    .io_d_out_15_valid_b(array_20_io_d_out_15_valid_b),
    .io_d_out_16_a(array_20_io_d_out_16_a),
    .io_d_out_16_valid_a(array_20_io_d_out_16_valid_a),
    .io_d_out_16_b(array_20_io_d_out_16_b),
    .io_d_out_16_valid_b(array_20_io_d_out_16_valid_b),
    .io_d_out_17_a(array_20_io_d_out_17_a),
    .io_d_out_17_valid_a(array_20_io_d_out_17_valid_a),
    .io_d_out_17_b(array_20_io_d_out_17_b),
    .io_d_out_17_valid_b(array_20_io_d_out_17_valid_b),
    .io_d_out_18_a(array_20_io_d_out_18_a),
    .io_d_out_18_valid_a(array_20_io_d_out_18_valid_a),
    .io_d_out_18_b(array_20_io_d_out_18_b),
    .io_d_out_18_valid_b(array_20_io_d_out_18_valid_b),
    .io_d_out_19_a(array_20_io_d_out_19_a),
    .io_d_out_19_valid_a(array_20_io_d_out_19_valid_a),
    .io_d_out_19_b(array_20_io_d_out_19_b),
    .io_d_out_19_valid_b(array_20_io_d_out_19_valid_b),
    .io_d_out_20_a(array_20_io_d_out_20_a),
    .io_d_out_20_valid_a(array_20_io_d_out_20_valid_a),
    .io_d_out_20_b(array_20_io_d_out_20_b),
    .io_d_out_20_valid_b(array_20_io_d_out_20_valid_b),
    .io_d_out_21_a(array_20_io_d_out_21_a),
    .io_d_out_21_valid_a(array_20_io_d_out_21_valid_a),
    .io_d_out_21_b(array_20_io_d_out_21_b),
    .io_d_out_21_valid_b(array_20_io_d_out_21_valid_b),
    .io_d_out_22_a(array_20_io_d_out_22_a),
    .io_d_out_22_valid_a(array_20_io_d_out_22_valid_a),
    .io_d_out_22_b(array_20_io_d_out_22_b),
    .io_d_out_22_valid_b(array_20_io_d_out_22_valid_b),
    .io_d_out_23_a(array_20_io_d_out_23_a),
    .io_d_out_23_valid_a(array_20_io_d_out_23_valid_a),
    .io_d_out_23_b(array_20_io_d_out_23_b),
    .io_d_out_23_valid_b(array_20_io_d_out_23_valid_b),
    .io_d_out_24_a(array_20_io_d_out_24_a),
    .io_d_out_24_valid_a(array_20_io_d_out_24_valid_a),
    .io_d_out_24_b(array_20_io_d_out_24_b),
    .io_d_out_24_valid_b(array_20_io_d_out_24_valid_b),
    .io_d_out_25_a(array_20_io_d_out_25_a),
    .io_d_out_25_valid_a(array_20_io_d_out_25_valid_a),
    .io_d_out_25_b(array_20_io_d_out_25_b),
    .io_d_out_25_valid_b(array_20_io_d_out_25_valid_b),
    .io_d_out_26_a(array_20_io_d_out_26_a),
    .io_d_out_26_valid_a(array_20_io_d_out_26_valid_a),
    .io_d_out_26_b(array_20_io_d_out_26_b),
    .io_d_out_26_valid_b(array_20_io_d_out_26_valid_b),
    .io_d_out_27_a(array_20_io_d_out_27_a),
    .io_d_out_27_valid_a(array_20_io_d_out_27_valid_a),
    .io_d_out_27_b(array_20_io_d_out_27_b),
    .io_d_out_27_valid_b(array_20_io_d_out_27_valid_b),
    .io_d_out_28_a(array_20_io_d_out_28_a),
    .io_d_out_28_valid_a(array_20_io_d_out_28_valid_a),
    .io_d_out_28_b(array_20_io_d_out_28_b),
    .io_d_out_28_valid_b(array_20_io_d_out_28_valid_b),
    .io_d_out_29_a(array_20_io_d_out_29_a),
    .io_d_out_29_valid_a(array_20_io_d_out_29_valid_a),
    .io_d_out_29_b(array_20_io_d_out_29_b),
    .io_d_out_29_valid_b(array_20_io_d_out_29_valid_b),
    .io_d_out_30_a(array_20_io_d_out_30_a),
    .io_d_out_30_valid_a(array_20_io_d_out_30_valid_a),
    .io_d_out_30_b(array_20_io_d_out_30_b),
    .io_d_out_30_valid_b(array_20_io_d_out_30_valid_b),
    .io_d_out_31_a(array_20_io_d_out_31_a),
    .io_d_out_31_valid_a(array_20_io_d_out_31_valid_a),
    .io_d_out_31_b(array_20_io_d_out_31_b),
    .io_d_out_31_valid_b(array_20_io_d_out_31_valid_b),
    .io_wr_en_mem1(array_20_io_wr_en_mem1),
    .io_wr_en_mem2(array_20_io_wr_en_mem2),
    .io_wr_en_mem3(array_20_io_wr_en_mem3),
    .io_wr_en_mem4(array_20_io_wr_en_mem4),
    .io_wr_en_mem5(array_20_io_wr_en_mem5),
    .io_wr_en_mem6(array_20_io_wr_en_mem6),
    .io_wr_instr_mem1(array_20_io_wr_instr_mem1),
    .io_wr_instr_mem2(array_20_io_wr_instr_mem2),
    .io_wr_instr_mem3(array_20_io_wr_instr_mem3),
    .io_wr_instr_mem4(array_20_io_wr_instr_mem4),
    .io_wr_instr_mem5(array_20_io_wr_instr_mem5),
    .io_wr_instr_mem6(array_20_io_wr_instr_mem6),
    .io_PC1_in(array_20_io_PC1_in),
    .io_PC6_out(array_20_io_PC6_out),
    .io_Addr_in(array_20_io_Addr_in),
    .io_Addr_out(array_20_io_Addr_out)
  );
  assign inputDataBuffer_0_validBit_MPORT_3_addr = inputDataBuffer_0_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_0_validBit_MPORT_3_data = inputDataBuffer_0_validBit[inputDataBuffer_0_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_0_validBit_MPORT_data = io_wr_D_inBuf_0_validBit;
  assign inputDataBuffer_0_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_0_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_0_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_0_data_MPORT_3_addr = inputDataBuffer_0_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_0_data_MPORT_3_data = inputDataBuffer_0_data[inputDataBuffer_0_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_0_data_MPORT_data = io_wr_D_inBuf_0_data;
  assign inputDataBuffer_0_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_0_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_0_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_1_validBit_MPORT_3_addr = inputDataBuffer_1_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_1_validBit_MPORT_3_data = inputDataBuffer_1_validBit[inputDataBuffer_1_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_1_validBit_MPORT_data = io_wr_D_inBuf_1_validBit;
  assign inputDataBuffer_1_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_1_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_1_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_1_data_MPORT_3_addr = inputDataBuffer_1_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_1_data_MPORT_3_data = inputDataBuffer_1_data[inputDataBuffer_1_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_1_data_MPORT_data = io_wr_D_inBuf_1_data;
  assign inputDataBuffer_1_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_1_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_1_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_2_validBit_MPORT_3_addr = inputDataBuffer_2_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_2_validBit_MPORT_3_data = inputDataBuffer_2_validBit[inputDataBuffer_2_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_2_validBit_MPORT_data = io_wr_D_inBuf_2_validBit;
  assign inputDataBuffer_2_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_2_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_2_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_2_data_MPORT_3_addr = inputDataBuffer_2_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_2_data_MPORT_3_data = inputDataBuffer_2_data[inputDataBuffer_2_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_2_data_MPORT_data = io_wr_D_inBuf_2_data;
  assign inputDataBuffer_2_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_2_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_2_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_3_validBit_MPORT_3_addr = inputDataBuffer_3_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_3_validBit_MPORT_3_data = inputDataBuffer_3_validBit[inputDataBuffer_3_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_3_validBit_MPORT_data = io_wr_D_inBuf_3_validBit;
  assign inputDataBuffer_3_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_3_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_3_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_3_data_MPORT_3_addr = inputDataBuffer_3_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_3_data_MPORT_3_data = inputDataBuffer_3_data[inputDataBuffer_3_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_3_data_MPORT_data = io_wr_D_inBuf_3_data;
  assign inputDataBuffer_3_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_3_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_3_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_4_validBit_MPORT_3_addr = inputDataBuffer_4_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_4_validBit_MPORT_3_data = inputDataBuffer_4_validBit[inputDataBuffer_4_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_4_validBit_MPORT_data = io_wr_D_inBuf_4_validBit;
  assign inputDataBuffer_4_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_4_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_4_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_4_data_MPORT_3_addr = inputDataBuffer_4_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_4_data_MPORT_3_data = inputDataBuffer_4_data[inputDataBuffer_4_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_4_data_MPORT_data = io_wr_D_inBuf_4_data;
  assign inputDataBuffer_4_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_4_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_4_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_5_validBit_MPORT_3_addr = inputDataBuffer_5_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_5_validBit_MPORT_3_data = inputDataBuffer_5_validBit[inputDataBuffer_5_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_5_validBit_MPORT_data = io_wr_D_inBuf_5_validBit;
  assign inputDataBuffer_5_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_5_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_5_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_5_data_MPORT_3_addr = inputDataBuffer_5_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_5_data_MPORT_3_data = inputDataBuffer_5_data[inputDataBuffer_5_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_5_data_MPORT_data = io_wr_D_inBuf_5_data;
  assign inputDataBuffer_5_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_5_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_5_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_6_validBit_MPORT_3_addr = inputDataBuffer_6_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_6_validBit_MPORT_3_data = inputDataBuffer_6_validBit[inputDataBuffer_6_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_6_validBit_MPORT_data = io_wr_D_inBuf_6_validBit;
  assign inputDataBuffer_6_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_6_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_6_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_6_data_MPORT_3_addr = inputDataBuffer_6_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_6_data_MPORT_3_data = inputDataBuffer_6_data[inputDataBuffer_6_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_6_data_MPORT_data = io_wr_D_inBuf_6_data;
  assign inputDataBuffer_6_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_6_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_6_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_7_validBit_MPORT_3_addr = inputDataBuffer_7_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_7_validBit_MPORT_3_data = inputDataBuffer_7_validBit[inputDataBuffer_7_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_7_validBit_MPORT_data = io_wr_D_inBuf_7_validBit;
  assign inputDataBuffer_7_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_7_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_7_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_7_data_MPORT_3_addr = inputDataBuffer_7_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_7_data_MPORT_3_data = inputDataBuffer_7_data[inputDataBuffer_7_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_7_data_MPORT_data = io_wr_D_inBuf_7_data;
  assign inputDataBuffer_7_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_7_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_7_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_8_validBit_MPORT_3_addr = inputDataBuffer_8_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_8_validBit_MPORT_3_data = inputDataBuffer_8_validBit[inputDataBuffer_8_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_8_validBit_MPORT_data = io_wr_D_inBuf_8_validBit;
  assign inputDataBuffer_8_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_8_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_8_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_8_data_MPORT_3_addr = inputDataBuffer_8_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_8_data_MPORT_3_data = inputDataBuffer_8_data[inputDataBuffer_8_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_8_data_MPORT_data = io_wr_D_inBuf_8_data;
  assign inputDataBuffer_8_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_8_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_8_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_9_validBit_MPORT_3_addr = inputDataBuffer_9_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_9_validBit_MPORT_3_data = inputDataBuffer_9_validBit[inputDataBuffer_9_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_9_validBit_MPORT_data = io_wr_D_inBuf_9_validBit;
  assign inputDataBuffer_9_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_9_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_9_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_9_data_MPORT_3_addr = inputDataBuffer_9_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_9_data_MPORT_3_data = inputDataBuffer_9_data[inputDataBuffer_9_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_9_data_MPORT_data = io_wr_D_inBuf_9_data;
  assign inputDataBuffer_9_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_9_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_9_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_10_validBit_MPORT_3_addr = inputDataBuffer_10_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_10_validBit_MPORT_3_data =
    inputDataBuffer_10_validBit[inputDataBuffer_10_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_10_validBit_MPORT_data = io_wr_D_inBuf_10_validBit;
  assign inputDataBuffer_10_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_10_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_10_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_10_data_MPORT_3_addr = inputDataBuffer_10_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_10_data_MPORT_3_data = inputDataBuffer_10_data[inputDataBuffer_10_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_10_data_MPORT_data = io_wr_D_inBuf_10_data;
  assign inputDataBuffer_10_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_10_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_10_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_11_validBit_MPORT_3_addr = inputDataBuffer_11_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_11_validBit_MPORT_3_data =
    inputDataBuffer_11_validBit[inputDataBuffer_11_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_11_validBit_MPORT_data = io_wr_D_inBuf_11_validBit;
  assign inputDataBuffer_11_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_11_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_11_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_11_data_MPORT_3_addr = inputDataBuffer_11_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_11_data_MPORT_3_data = inputDataBuffer_11_data[inputDataBuffer_11_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_11_data_MPORT_data = io_wr_D_inBuf_11_data;
  assign inputDataBuffer_11_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_11_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_11_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_12_validBit_MPORT_3_addr = inputDataBuffer_12_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_12_validBit_MPORT_3_data =
    inputDataBuffer_12_validBit[inputDataBuffer_12_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_12_validBit_MPORT_data = io_wr_D_inBuf_12_validBit;
  assign inputDataBuffer_12_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_12_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_12_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_12_data_MPORT_3_addr = inputDataBuffer_12_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_12_data_MPORT_3_data = inputDataBuffer_12_data[inputDataBuffer_12_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_12_data_MPORT_data = io_wr_D_inBuf_12_data;
  assign inputDataBuffer_12_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_12_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_12_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_13_validBit_MPORT_3_addr = inputDataBuffer_13_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_13_validBit_MPORT_3_data =
    inputDataBuffer_13_validBit[inputDataBuffer_13_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_13_validBit_MPORT_data = io_wr_D_inBuf_13_validBit;
  assign inputDataBuffer_13_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_13_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_13_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_13_data_MPORT_3_addr = inputDataBuffer_13_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_13_data_MPORT_3_data = inputDataBuffer_13_data[inputDataBuffer_13_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_13_data_MPORT_data = io_wr_D_inBuf_13_data;
  assign inputDataBuffer_13_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_13_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_13_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_14_validBit_MPORT_3_addr = inputDataBuffer_14_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_14_validBit_MPORT_3_data =
    inputDataBuffer_14_validBit[inputDataBuffer_14_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_14_validBit_MPORT_data = io_wr_D_inBuf_14_validBit;
  assign inputDataBuffer_14_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_14_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_14_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_14_data_MPORT_3_addr = inputDataBuffer_14_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_14_data_MPORT_3_data = inputDataBuffer_14_data[inputDataBuffer_14_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_14_data_MPORT_data = io_wr_D_inBuf_14_data;
  assign inputDataBuffer_14_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_14_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_14_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_15_validBit_MPORT_3_addr = inputDataBuffer_15_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_15_validBit_MPORT_3_data =
    inputDataBuffer_15_validBit[inputDataBuffer_15_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_15_validBit_MPORT_data = io_wr_D_inBuf_15_validBit;
  assign inputDataBuffer_15_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_15_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_15_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_15_data_MPORT_3_addr = inputDataBuffer_15_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_15_data_MPORT_3_data = inputDataBuffer_15_data[inputDataBuffer_15_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_15_data_MPORT_data = io_wr_D_inBuf_15_data;
  assign inputDataBuffer_15_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_15_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_15_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_16_validBit_MPORT_3_addr = inputDataBuffer_16_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_16_validBit_MPORT_3_data =
    inputDataBuffer_16_validBit[inputDataBuffer_16_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_16_validBit_MPORT_data = io_wr_D_inBuf_16_validBit;
  assign inputDataBuffer_16_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_16_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_16_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_16_data_MPORT_3_addr = inputDataBuffer_16_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_16_data_MPORT_3_data = inputDataBuffer_16_data[inputDataBuffer_16_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_16_data_MPORT_data = io_wr_D_inBuf_16_data;
  assign inputDataBuffer_16_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_16_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_16_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_17_validBit_MPORT_3_addr = inputDataBuffer_17_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_17_validBit_MPORT_3_data =
    inputDataBuffer_17_validBit[inputDataBuffer_17_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_17_validBit_MPORT_data = io_wr_D_inBuf_17_validBit;
  assign inputDataBuffer_17_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_17_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_17_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_17_data_MPORT_3_addr = inputDataBuffer_17_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_17_data_MPORT_3_data = inputDataBuffer_17_data[inputDataBuffer_17_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_17_data_MPORT_data = io_wr_D_inBuf_17_data;
  assign inputDataBuffer_17_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_17_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_17_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_18_validBit_MPORT_3_addr = inputDataBuffer_18_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_18_validBit_MPORT_3_data =
    inputDataBuffer_18_validBit[inputDataBuffer_18_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_18_validBit_MPORT_data = io_wr_D_inBuf_18_validBit;
  assign inputDataBuffer_18_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_18_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_18_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_18_data_MPORT_3_addr = inputDataBuffer_18_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_18_data_MPORT_3_data = inputDataBuffer_18_data[inputDataBuffer_18_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_18_data_MPORT_data = io_wr_D_inBuf_18_data;
  assign inputDataBuffer_18_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_18_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_18_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_19_validBit_MPORT_3_addr = inputDataBuffer_19_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_19_validBit_MPORT_3_data =
    inputDataBuffer_19_validBit[inputDataBuffer_19_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_19_validBit_MPORT_data = io_wr_D_inBuf_19_validBit;
  assign inputDataBuffer_19_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_19_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_19_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_19_data_MPORT_3_addr = inputDataBuffer_19_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_19_data_MPORT_3_data = inputDataBuffer_19_data[inputDataBuffer_19_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_19_data_MPORT_data = io_wr_D_inBuf_19_data;
  assign inputDataBuffer_19_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_19_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_19_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_20_validBit_MPORT_3_addr = inputDataBuffer_20_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_20_validBit_MPORT_3_data =
    inputDataBuffer_20_validBit[inputDataBuffer_20_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_20_validBit_MPORT_data = io_wr_D_inBuf_20_validBit;
  assign inputDataBuffer_20_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_20_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_20_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_20_data_MPORT_3_addr = inputDataBuffer_20_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_20_data_MPORT_3_data = inputDataBuffer_20_data[inputDataBuffer_20_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_20_data_MPORT_data = io_wr_D_inBuf_20_data;
  assign inputDataBuffer_20_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_20_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_20_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_21_validBit_MPORT_3_addr = inputDataBuffer_21_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_21_validBit_MPORT_3_data =
    inputDataBuffer_21_validBit[inputDataBuffer_21_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_21_validBit_MPORT_data = io_wr_D_inBuf_21_validBit;
  assign inputDataBuffer_21_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_21_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_21_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_21_data_MPORT_3_addr = inputDataBuffer_21_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_21_data_MPORT_3_data = inputDataBuffer_21_data[inputDataBuffer_21_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_21_data_MPORT_data = io_wr_D_inBuf_21_data;
  assign inputDataBuffer_21_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_21_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_21_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_22_validBit_MPORT_3_addr = inputDataBuffer_22_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_22_validBit_MPORT_3_data =
    inputDataBuffer_22_validBit[inputDataBuffer_22_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_22_validBit_MPORT_data = io_wr_D_inBuf_22_validBit;
  assign inputDataBuffer_22_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_22_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_22_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_22_data_MPORT_3_addr = inputDataBuffer_22_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_22_data_MPORT_3_data = inputDataBuffer_22_data[inputDataBuffer_22_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_22_data_MPORT_data = io_wr_D_inBuf_22_data;
  assign inputDataBuffer_22_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_22_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_22_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_23_validBit_MPORT_3_addr = inputDataBuffer_23_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_23_validBit_MPORT_3_data =
    inputDataBuffer_23_validBit[inputDataBuffer_23_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_23_validBit_MPORT_data = io_wr_D_inBuf_23_validBit;
  assign inputDataBuffer_23_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_23_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_23_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_23_data_MPORT_3_addr = inputDataBuffer_23_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_23_data_MPORT_3_data = inputDataBuffer_23_data[inputDataBuffer_23_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_23_data_MPORT_data = io_wr_D_inBuf_23_data;
  assign inputDataBuffer_23_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_23_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_23_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_24_validBit_MPORT_3_addr = inputDataBuffer_24_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_24_validBit_MPORT_3_data =
    inputDataBuffer_24_validBit[inputDataBuffer_24_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_24_validBit_MPORT_data = io_wr_D_inBuf_24_validBit;
  assign inputDataBuffer_24_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_24_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_24_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_24_data_MPORT_3_addr = inputDataBuffer_24_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_24_data_MPORT_3_data = inputDataBuffer_24_data[inputDataBuffer_24_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_24_data_MPORT_data = io_wr_D_inBuf_24_data;
  assign inputDataBuffer_24_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_24_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_24_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_25_validBit_MPORT_3_addr = inputDataBuffer_25_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_25_validBit_MPORT_3_data =
    inputDataBuffer_25_validBit[inputDataBuffer_25_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_25_validBit_MPORT_data = io_wr_D_inBuf_25_validBit;
  assign inputDataBuffer_25_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_25_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_25_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_25_data_MPORT_3_addr = inputDataBuffer_25_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_25_data_MPORT_3_data = inputDataBuffer_25_data[inputDataBuffer_25_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_25_data_MPORT_data = io_wr_D_inBuf_25_data;
  assign inputDataBuffer_25_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_25_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_25_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_26_validBit_MPORT_3_addr = inputDataBuffer_26_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_26_validBit_MPORT_3_data =
    inputDataBuffer_26_validBit[inputDataBuffer_26_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_26_validBit_MPORT_data = io_wr_D_inBuf_26_validBit;
  assign inputDataBuffer_26_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_26_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_26_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_26_data_MPORT_3_addr = inputDataBuffer_26_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_26_data_MPORT_3_data = inputDataBuffer_26_data[inputDataBuffer_26_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_26_data_MPORT_data = io_wr_D_inBuf_26_data;
  assign inputDataBuffer_26_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_26_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_26_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_27_validBit_MPORT_3_addr = inputDataBuffer_27_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_27_validBit_MPORT_3_data =
    inputDataBuffer_27_validBit[inputDataBuffer_27_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_27_validBit_MPORT_data = io_wr_D_inBuf_27_validBit;
  assign inputDataBuffer_27_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_27_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_27_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_27_data_MPORT_3_addr = inputDataBuffer_27_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_27_data_MPORT_3_data = inputDataBuffer_27_data[inputDataBuffer_27_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_27_data_MPORT_data = io_wr_D_inBuf_27_data;
  assign inputDataBuffer_27_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_27_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_27_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_28_validBit_MPORT_3_addr = inputDataBuffer_28_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_28_validBit_MPORT_3_data =
    inputDataBuffer_28_validBit[inputDataBuffer_28_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_28_validBit_MPORT_data = io_wr_D_inBuf_28_validBit;
  assign inputDataBuffer_28_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_28_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_28_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_28_data_MPORT_3_addr = inputDataBuffer_28_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_28_data_MPORT_3_data = inputDataBuffer_28_data[inputDataBuffer_28_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_28_data_MPORT_data = io_wr_D_inBuf_28_data;
  assign inputDataBuffer_28_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_28_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_28_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_29_validBit_MPORT_3_addr = inputDataBuffer_29_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_29_validBit_MPORT_3_data =
    inputDataBuffer_29_validBit[inputDataBuffer_29_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_29_validBit_MPORT_data = io_wr_D_inBuf_29_validBit;
  assign inputDataBuffer_29_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_29_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_29_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_29_data_MPORT_3_addr = inputDataBuffer_29_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_29_data_MPORT_3_data = inputDataBuffer_29_data[inputDataBuffer_29_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_29_data_MPORT_data = io_wr_D_inBuf_29_data;
  assign inputDataBuffer_29_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_29_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_29_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_30_validBit_MPORT_3_addr = inputDataBuffer_30_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_30_validBit_MPORT_3_data =
    inputDataBuffer_30_validBit[inputDataBuffer_30_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_30_validBit_MPORT_data = io_wr_D_inBuf_30_validBit;
  assign inputDataBuffer_30_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_30_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_30_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_30_data_MPORT_3_addr = inputDataBuffer_30_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_30_data_MPORT_3_data = inputDataBuffer_30_data[inputDataBuffer_30_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_30_data_MPORT_data = io_wr_D_inBuf_30_data;
  assign inputDataBuffer_30_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_30_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_30_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_31_validBit_MPORT_3_addr = inputDataBuffer_31_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_31_validBit_MPORT_3_data =
    inputDataBuffer_31_validBit[inputDataBuffer_31_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_31_validBit_MPORT_data = io_wr_D_inBuf_31_validBit;
  assign inputDataBuffer_31_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_31_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_31_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_31_data_MPORT_3_addr = inputDataBuffer_31_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_31_data_MPORT_3_data = inputDataBuffer_31_data[inputDataBuffer_31_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_31_data_MPORT_data = io_wr_D_inBuf_31_data;
  assign inputDataBuffer_31_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_31_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_31_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_32_validBit_MPORT_3_addr = inputDataBuffer_32_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_32_validBit_MPORT_3_data =
    inputDataBuffer_32_validBit[inputDataBuffer_32_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_32_validBit_MPORT_data = io_wr_D_inBuf_32_validBit;
  assign inputDataBuffer_32_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_32_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_32_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_32_data_MPORT_3_addr = inputDataBuffer_32_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_32_data_MPORT_3_data = inputDataBuffer_32_data[inputDataBuffer_32_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_32_data_MPORT_data = io_wr_D_inBuf_32_data;
  assign inputDataBuffer_32_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_32_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_32_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_33_validBit_MPORT_3_addr = inputDataBuffer_33_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_33_validBit_MPORT_3_data =
    inputDataBuffer_33_validBit[inputDataBuffer_33_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_33_validBit_MPORT_data = io_wr_D_inBuf_33_validBit;
  assign inputDataBuffer_33_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_33_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_33_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_33_data_MPORT_3_addr = inputDataBuffer_33_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_33_data_MPORT_3_data = inputDataBuffer_33_data[inputDataBuffer_33_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_33_data_MPORT_data = io_wr_D_inBuf_33_data;
  assign inputDataBuffer_33_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_33_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_33_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_34_validBit_MPORT_3_addr = inputDataBuffer_34_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_34_validBit_MPORT_3_data =
    inputDataBuffer_34_validBit[inputDataBuffer_34_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_34_validBit_MPORT_data = io_wr_D_inBuf_34_validBit;
  assign inputDataBuffer_34_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_34_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_34_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_34_data_MPORT_3_addr = inputDataBuffer_34_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_34_data_MPORT_3_data = inputDataBuffer_34_data[inputDataBuffer_34_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_34_data_MPORT_data = io_wr_D_inBuf_34_data;
  assign inputDataBuffer_34_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_34_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_34_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_35_validBit_MPORT_3_addr = inputDataBuffer_35_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_35_validBit_MPORT_3_data =
    inputDataBuffer_35_validBit[inputDataBuffer_35_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_35_validBit_MPORT_data = io_wr_D_inBuf_35_validBit;
  assign inputDataBuffer_35_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_35_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_35_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_35_data_MPORT_3_addr = inputDataBuffer_35_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_35_data_MPORT_3_data = inputDataBuffer_35_data[inputDataBuffer_35_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_35_data_MPORT_data = io_wr_D_inBuf_35_data;
  assign inputDataBuffer_35_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_35_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_35_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_36_validBit_MPORT_3_addr = inputDataBuffer_36_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_36_validBit_MPORT_3_data =
    inputDataBuffer_36_validBit[inputDataBuffer_36_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_36_validBit_MPORT_data = io_wr_D_inBuf_36_validBit;
  assign inputDataBuffer_36_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_36_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_36_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_36_data_MPORT_3_addr = inputDataBuffer_36_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_36_data_MPORT_3_data = inputDataBuffer_36_data[inputDataBuffer_36_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_36_data_MPORT_data = io_wr_D_inBuf_36_data;
  assign inputDataBuffer_36_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_36_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_36_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_37_validBit_MPORT_3_addr = inputDataBuffer_37_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_37_validBit_MPORT_3_data =
    inputDataBuffer_37_validBit[inputDataBuffer_37_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_37_validBit_MPORT_data = io_wr_D_inBuf_37_validBit;
  assign inputDataBuffer_37_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_37_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_37_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_37_data_MPORT_3_addr = inputDataBuffer_37_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_37_data_MPORT_3_data = inputDataBuffer_37_data[inputDataBuffer_37_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_37_data_MPORT_data = io_wr_D_inBuf_37_data;
  assign inputDataBuffer_37_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_37_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_37_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_38_validBit_MPORT_3_addr = inputDataBuffer_38_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_38_validBit_MPORT_3_data =
    inputDataBuffer_38_validBit[inputDataBuffer_38_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_38_validBit_MPORT_data = io_wr_D_inBuf_38_validBit;
  assign inputDataBuffer_38_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_38_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_38_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_38_data_MPORT_3_addr = inputDataBuffer_38_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_38_data_MPORT_3_data = inputDataBuffer_38_data[inputDataBuffer_38_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_38_data_MPORT_data = io_wr_D_inBuf_38_data;
  assign inputDataBuffer_38_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_38_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_38_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_39_validBit_MPORT_3_addr = inputDataBuffer_39_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_39_validBit_MPORT_3_data =
    inputDataBuffer_39_validBit[inputDataBuffer_39_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_39_validBit_MPORT_data = io_wr_D_inBuf_39_validBit;
  assign inputDataBuffer_39_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_39_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_39_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_39_data_MPORT_3_addr = inputDataBuffer_39_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_39_data_MPORT_3_data = inputDataBuffer_39_data[inputDataBuffer_39_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_39_data_MPORT_data = io_wr_D_inBuf_39_data;
  assign inputDataBuffer_39_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_39_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_39_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_40_validBit_MPORT_3_addr = inputDataBuffer_40_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_40_validBit_MPORT_3_data =
    inputDataBuffer_40_validBit[inputDataBuffer_40_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_40_validBit_MPORT_data = io_wr_D_inBuf_40_validBit;
  assign inputDataBuffer_40_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_40_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_40_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_40_data_MPORT_3_addr = inputDataBuffer_40_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_40_data_MPORT_3_data = inputDataBuffer_40_data[inputDataBuffer_40_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_40_data_MPORT_data = io_wr_D_inBuf_40_data;
  assign inputDataBuffer_40_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_40_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_40_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_41_validBit_MPORT_3_addr = inputDataBuffer_41_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_41_validBit_MPORT_3_data =
    inputDataBuffer_41_validBit[inputDataBuffer_41_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_41_validBit_MPORT_data = io_wr_D_inBuf_41_validBit;
  assign inputDataBuffer_41_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_41_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_41_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_41_data_MPORT_3_addr = inputDataBuffer_41_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_41_data_MPORT_3_data = inputDataBuffer_41_data[inputDataBuffer_41_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_41_data_MPORT_data = io_wr_D_inBuf_41_data;
  assign inputDataBuffer_41_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_41_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_41_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_42_validBit_MPORT_3_addr = inputDataBuffer_42_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_42_validBit_MPORT_3_data =
    inputDataBuffer_42_validBit[inputDataBuffer_42_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_42_validBit_MPORT_data = io_wr_D_inBuf_42_validBit;
  assign inputDataBuffer_42_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_42_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_42_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_42_data_MPORT_3_addr = inputDataBuffer_42_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_42_data_MPORT_3_data = inputDataBuffer_42_data[inputDataBuffer_42_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_42_data_MPORT_data = io_wr_D_inBuf_42_data;
  assign inputDataBuffer_42_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_42_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_42_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_43_validBit_MPORT_3_addr = inputDataBuffer_43_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_43_validBit_MPORT_3_data =
    inputDataBuffer_43_validBit[inputDataBuffer_43_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_43_validBit_MPORT_data = io_wr_D_inBuf_43_validBit;
  assign inputDataBuffer_43_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_43_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_43_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_43_data_MPORT_3_addr = inputDataBuffer_43_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_43_data_MPORT_3_data = inputDataBuffer_43_data[inputDataBuffer_43_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_43_data_MPORT_data = io_wr_D_inBuf_43_data;
  assign inputDataBuffer_43_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_43_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_43_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_44_validBit_MPORT_3_addr = inputDataBuffer_44_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_44_validBit_MPORT_3_data =
    inputDataBuffer_44_validBit[inputDataBuffer_44_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_44_validBit_MPORT_data = io_wr_D_inBuf_44_validBit;
  assign inputDataBuffer_44_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_44_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_44_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_44_data_MPORT_3_addr = inputDataBuffer_44_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_44_data_MPORT_3_data = inputDataBuffer_44_data[inputDataBuffer_44_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_44_data_MPORT_data = io_wr_D_inBuf_44_data;
  assign inputDataBuffer_44_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_44_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_44_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_45_validBit_MPORT_3_addr = inputDataBuffer_45_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_45_validBit_MPORT_3_data =
    inputDataBuffer_45_validBit[inputDataBuffer_45_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_45_validBit_MPORT_data = io_wr_D_inBuf_45_validBit;
  assign inputDataBuffer_45_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_45_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_45_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_45_data_MPORT_3_addr = inputDataBuffer_45_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_45_data_MPORT_3_data = inputDataBuffer_45_data[inputDataBuffer_45_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_45_data_MPORT_data = io_wr_D_inBuf_45_data;
  assign inputDataBuffer_45_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_45_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_45_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_46_validBit_MPORT_3_addr = inputDataBuffer_46_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_46_validBit_MPORT_3_data =
    inputDataBuffer_46_validBit[inputDataBuffer_46_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_46_validBit_MPORT_data = io_wr_D_inBuf_46_validBit;
  assign inputDataBuffer_46_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_46_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_46_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_46_data_MPORT_3_addr = inputDataBuffer_46_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_46_data_MPORT_3_data = inputDataBuffer_46_data[inputDataBuffer_46_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_46_data_MPORT_data = io_wr_D_inBuf_46_data;
  assign inputDataBuffer_46_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_46_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_46_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_47_validBit_MPORT_3_addr = inputDataBuffer_47_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_47_validBit_MPORT_3_data =
    inputDataBuffer_47_validBit[inputDataBuffer_47_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_47_validBit_MPORT_data = io_wr_D_inBuf_47_validBit;
  assign inputDataBuffer_47_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_47_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_47_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_47_data_MPORT_3_addr = inputDataBuffer_47_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_47_data_MPORT_3_data = inputDataBuffer_47_data[inputDataBuffer_47_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_47_data_MPORT_data = io_wr_D_inBuf_47_data;
  assign inputDataBuffer_47_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_47_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_47_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_48_validBit_MPORT_3_addr = inputDataBuffer_48_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_48_validBit_MPORT_3_data =
    inputDataBuffer_48_validBit[inputDataBuffer_48_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_48_validBit_MPORT_data = io_wr_D_inBuf_48_validBit;
  assign inputDataBuffer_48_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_48_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_48_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_48_data_MPORT_3_addr = inputDataBuffer_48_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_48_data_MPORT_3_data = inputDataBuffer_48_data[inputDataBuffer_48_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_48_data_MPORT_data = io_wr_D_inBuf_48_data;
  assign inputDataBuffer_48_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_48_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_48_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_49_validBit_MPORT_3_addr = inputDataBuffer_49_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_49_validBit_MPORT_3_data =
    inputDataBuffer_49_validBit[inputDataBuffer_49_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_49_validBit_MPORT_data = io_wr_D_inBuf_49_validBit;
  assign inputDataBuffer_49_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_49_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_49_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_49_data_MPORT_3_addr = inputDataBuffer_49_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_49_data_MPORT_3_data = inputDataBuffer_49_data[inputDataBuffer_49_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_49_data_MPORT_data = io_wr_D_inBuf_49_data;
  assign inputDataBuffer_49_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_49_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_49_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_50_validBit_MPORT_3_addr = inputDataBuffer_50_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_50_validBit_MPORT_3_data =
    inputDataBuffer_50_validBit[inputDataBuffer_50_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_50_validBit_MPORT_data = io_wr_D_inBuf_50_validBit;
  assign inputDataBuffer_50_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_50_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_50_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_50_data_MPORT_3_addr = inputDataBuffer_50_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_50_data_MPORT_3_data = inputDataBuffer_50_data[inputDataBuffer_50_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_50_data_MPORT_data = io_wr_D_inBuf_50_data;
  assign inputDataBuffer_50_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_50_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_50_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_51_validBit_MPORT_3_addr = inputDataBuffer_51_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_51_validBit_MPORT_3_data =
    inputDataBuffer_51_validBit[inputDataBuffer_51_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_51_validBit_MPORT_data = io_wr_D_inBuf_51_validBit;
  assign inputDataBuffer_51_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_51_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_51_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_51_data_MPORT_3_addr = inputDataBuffer_51_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_51_data_MPORT_3_data = inputDataBuffer_51_data[inputDataBuffer_51_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_51_data_MPORT_data = io_wr_D_inBuf_51_data;
  assign inputDataBuffer_51_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_51_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_51_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_52_validBit_MPORT_3_addr = inputDataBuffer_52_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_52_validBit_MPORT_3_data =
    inputDataBuffer_52_validBit[inputDataBuffer_52_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_52_validBit_MPORT_data = io_wr_D_inBuf_52_validBit;
  assign inputDataBuffer_52_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_52_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_52_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_52_data_MPORT_3_addr = inputDataBuffer_52_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_52_data_MPORT_3_data = inputDataBuffer_52_data[inputDataBuffer_52_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_52_data_MPORT_data = io_wr_D_inBuf_52_data;
  assign inputDataBuffer_52_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_52_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_52_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_53_validBit_MPORT_3_addr = inputDataBuffer_53_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_53_validBit_MPORT_3_data =
    inputDataBuffer_53_validBit[inputDataBuffer_53_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_53_validBit_MPORT_data = io_wr_D_inBuf_53_validBit;
  assign inputDataBuffer_53_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_53_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_53_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_53_data_MPORT_3_addr = inputDataBuffer_53_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_53_data_MPORT_3_data = inputDataBuffer_53_data[inputDataBuffer_53_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_53_data_MPORT_data = io_wr_D_inBuf_53_data;
  assign inputDataBuffer_53_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_53_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_53_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_54_validBit_MPORT_3_addr = inputDataBuffer_54_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_54_validBit_MPORT_3_data =
    inputDataBuffer_54_validBit[inputDataBuffer_54_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_54_validBit_MPORT_data = io_wr_D_inBuf_54_validBit;
  assign inputDataBuffer_54_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_54_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_54_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_54_data_MPORT_3_addr = inputDataBuffer_54_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_54_data_MPORT_3_data = inputDataBuffer_54_data[inputDataBuffer_54_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_54_data_MPORT_data = io_wr_D_inBuf_54_data;
  assign inputDataBuffer_54_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_54_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_54_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_55_validBit_MPORT_3_addr = inputDataBuffer_55_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_55_validBit_MPORT_3_data =
    inputDataBuffer_55_validBit[inputDataBuffer_55_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_55_validBit_MPORT_data = io_wr_D_inBuf_55_validBit;
  assign inputDataBuffer_55_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_55_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_55_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_55_data_MPORT_3_addr = inputDataBuffer_55_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_55_data_MPORT_3_data = inputDataBuffer_55_data[inputDataBuffer_55_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_55_data_MPORT_data = io_wr_D_inBuf_55_data;
  assign inputDataBuffer_55_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_55_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_55_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_56_validBit_MPORT_3_addr = inputDataBuffer_56_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_56_validBit_MPORT_3_data =
    inputDataBuffer_56_validBit[inputDataBuffer_56_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_56_validBit_MPORT_data = io_wr_D_inBuf_56_validBit;
  assign inputDataBuffer_56_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_56_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_56_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_56_data_MPORT_3_addr = inputDataBuffer_56_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_56_data_MPORT_3_data = inputDataBuffer_56_data[inputDataBuffer_56_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_56_data_MPORT_data = io_wr_D_inBuf_56_data;
  assign inputDataBuffer_56_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_56_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_56_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_57_validBit_MPORT_3_addr = inputDataBuffer_57_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_57_validBit_MPORT_3_data =
    inputDataBuffer_57_validBit[inputDataBuffer_57_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_57_validBit_MPORT_data = io_wr_D_inBuf_57_validBit;
  assign inputDataBuffer_57_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_57_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_57_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_57_data_MPORT_3_addr = inputDataBuffer_57_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_57_data_MPORT_3_data = inputDataBuffer_57_data[inputDataBuffer_57_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_57_data_MPORT_data = io_wr_D_inBuf_57_data;
  assign inputDataBuffer_57_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_57_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_57_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_58_validBit_MPORT_3_addr = inputDataBuffer_58_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_58_validBit_MPORT_3_data =
    inputDataBuffer_58_validBit[inputDataBuffer_58_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_58_validBit_MPORT_data = io_wr_D_inBuf_58_validBit;
  assign inputDataBuffer_58_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_58_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_58_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_58_data_MPORT_3_addr = inputDataBuffer_58_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_58_data_MPORT_3_data = inputDataBuffer_58_data[inputDataBuffer_58_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_58_data_MPORT_data = io_wr_D_inBuf_58_data;
  assign inputDataBuffer_58_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_58_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_58_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_59_validBit_MPORT_3_addr = inputDataBuffer_59_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_59_validBit_MPORT_3_data =
    inputDataBuffer_59_validBit[inputDataBuffer_59_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_59_validBit_MPORT_data = io_wr_D_inBuf_59_validBit;
  assign inputDataBuffer_59_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_59_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_59_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_59_data_MPORT_3_addr = inputDataBuffer_59_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_59_data_MPORT_3_data = inputDataBuffer_59_data[inputDataBuffer_59_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_59_data_MPORT_data = io_wr_D_inBuf_59_data;
  assign inputDataBuffer_59_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_59_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_59_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_60_validBit_MPORT_3_addr = inputDataBuffer_60_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_60_validBit_MPORT_3_data =
    inputDataBuffer_60_validBit[inputDataBuffer_60_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_60_validBit_MPORT_data = io_wr_D_inBuf_60_validBit;
  assign inputDataBuffer_60_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_60_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_60_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_60_data_MPORT_3_addr = inputDataBuffer_60_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_60_data_MPORT_3_data = inputDataBuffer_60_data[inputDataBuffer_60_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_60_data_MPORT_data = io_wr_D_inBuf_60_data;
  assign inputDataBuffer_60_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_60_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_60_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_61_validBit_MPORT_3_addr = inputDataBuffer_61_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_61_validBit_MPORT_3_data =
    inputDataBuffer_61_validBit[inputDataBuffer_61_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_61_validBit_MPORT_data = io_wr_D_inBuf_61_validBit;
  assign inputDataBuffer_61_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_61_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_61_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_61_data_MPORT_3_addr = inputDataBuffer_61_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_61_data_MPORT_3_data = inputDataBuffer_61_data[inputDataBuffer_61_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_61_data_MPORT_data = io_wr_D_inBuf_61_data;
  assign inputDataBuffer_61_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_61_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_61_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_62_validBit_MPORT_3_addr = inputDataBuffer_62_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_62_validBit_MPORT_3_data =
    inputDataBuffer_62_validBit[inputDataBuffer_62_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_62_validBit_MPORT_data = io_wr_D_inBuf_62_validBit;
  assign inputDataBuffer_62_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_62_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_62_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_62_data_MPORT_3_addr = inputDataBuffer_62_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_62_data_MPORT_3_data = inputDataBuffer_62_data[inputDataBuffer_62_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_62_data_MPORT_data = io_wr_D_inBuf_62_data;
  assign inputDataBuffer_62_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_62_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_62_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_63_validBit_MPORT_3_addr = inputDataBuffer_63_validBit_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_63_validBit_MPORT_3_data =
    inputDataBuffer_63_validBit[inputDataBuffer_63_validBit_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_63_validBit_MPORT_data = io_wr_D_inBuf_63_validBit;
  assign inputDataBuffer_63_validBit_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_63_validBit_MPORT_mask = 1'h1;
  assign inputDataBuffer_63_validBit_MPORT_en = io_wr_Addr_inBuf_en;
  assign inputDataBuffer_63_data_MPORT_3_addr = inputDataBuffer_63_data_MPORT_3_addr_pipe_0;
  assign inputDataBuffer_63_data_MPORT_3_data = inputDataBuffer_63_data[inputDataBuffer_63_data_MPORT_3_addr]; // @[BP.scala 42:36]
  assign inputDataBuffer_63_data_MPORT_data = io_wr_D_inBuf_63_data;
  assign inputDataBuffer_63_data_MPORT_addr = wr_Addr_inBuf;
  assign inputDataBuffer_63_data_MPORT_mask = 1'h1;
  assign inputDataBuffer_63_data_MPORT_en = io_wr_Addr_inBuf_en;
  assign outputDataBuffer_0_validBit_MPORT_2_addr = outputDataBuffer_0_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_0_validBit_MPORT_2_data =
    outputDataBuffer_0_validBit[outputDataBuffer_0_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_0_validBit_MPORT_4_data = wr_D_outBuf_0_validBit;
  assign outputDataBuffer_0_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_0_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_0_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_0_data_MPORT_2_addr = outputDataBuffer_0_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_0_data_MPORT_2_data = outputDataBuffer_0_data[outputDataBuffer_0_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_0_data_MPORT_4_data = wr_D_outBuf_0_data;
  assign outputDataBuffer_0_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_0_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_0_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_1_validBit_MPORT_2_addr = outputDataBuffer_1_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_1_validBit_MPORT_2_data =
    outputDataBuffer_1_validBit[outputDataBuffer_1_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_1_validBit_MPORT_4_data = wr_D_outBuf_1_validBit;
  assign outputDataBuffer_1_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_1_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_1_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_1_data_MPORT_2_addr = outputDataBuffer_1_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_1_data_MPORT_2_data = outputDataBuffer_1_data[outputDataBuffer_1_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_1_data_MPORT_4_data = wr_D_outBuf_1_data;
  assign outputDataBuffer_1_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_1_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_1_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_2_validBit_MPORT_2_addr = outputDataBuffer_2_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_2_validBit_MPORT_2_data =
    outputDataBuffer_2_validBit[outputDataBuffer_2_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_2_validBit_MPORT_4_data = wr_D_outBuf_2_validBit;
  assign outputDataBuffer_2_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_2_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_2_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_2_data_MPORT_2_addr = outputDataBuffer_2_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_2_data_MPORT_2_data = outputDataBuffer_2_data[outputDataBuffer_2_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_2_data_MPORT_4_data = wr_D_outBuf_2_data;
  assign outputDataBuffer_2_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_2_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_2_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_3_validBit_MPORT_2_addr = outputDataBuffer_3_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_3_validBit_MPORT_2_data =
    outputDataBuffer_3_validBit[outputDataBuffer_3_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_3_validBit_MPORT_4_data = wr_D_outBuf_3_validBit;
  assign outputDataBuffer_3_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_3_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_3_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_3_data_MPORT_2_addr = outputDataBuffer_3_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_3_data_MPORT_2_data = outputDataBuffer_3_data[outputDataBuffer_3_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_3_data_MPORT_4_data = wr_D_outBuf_3_data;
  assign outputDataBuffer_3_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_3_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_3_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_4_validBit_MPORT_2_addr = outputDataBuffer_4_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_4_validBit_MPORT_2_data =
    outputDataBuffer_4_validBit[outputDataBuffer_4_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_4_validBit_MPORT_4_data = wr_D_outBuf_4_validBit;
  assign outputDataBuffer_4_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_4_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_4_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_4_data_MPORT_2_addr = outputDataBuffer_4_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_4_data_MPORT_2_data = outputDataBuffer_4_data[outputDataBuffer_4_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_4_data_MPORT_4_data = wr_D_outBuf_4_data;
  assign outputDataBuffer_4_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_4_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_4_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_5_validBit_MPORT_2_addr = outputDataBuffer_5_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_5_validBit_MPORT_2_data =
    outputDataBuffer_5_validBit[outputDataBuffer_5_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_5_validBit_MPORT_4_data = wr_D_outBuf_5_validBit;
  assign outputDataBuffer_5_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_5_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_5_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_5_data_MPORT_2_addr = outputDataBuffer_5_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_5_data_MPORT_2_data = outputDataBuffer_5_data[outputDataBuffer_5_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_5_data_MPORT_4_data = wr_D_outBuf_5_data;
  assign outputDataBuffer_5_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_5_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_5_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_6_validBit_MPORT_2_addr = outputDataBuffer_6_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_6_validBit_MPORT_2_data =
    outputDataBuffer_6_validBit[outputDataBuffer_6_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_6_validBit_MPORT_4_data = wr_D_outBuf_6_validBit;
  assign outputDataBuffer_6_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_6_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_6_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_6_data_MPORT_2_addr = outputDataBuffer_6_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_6_data_MPORT_2_data = outputDataBuffer_6_data[outputDataBuffer_6_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_6_data_MPORT_4_data = wr_D_outBuf_6_data;
  assign outputDataBuffer_6_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_6_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_6_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_7_validBit_MPORT_2_addr = outputDataBuffer_7_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_7_validBit_MPORT_2_data =
    outputDataBuffer_7_validBit[outputDataBuffer_7_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_7_validBit_MPORT_4_data = wr_D_outBuf_7_validBit;
  assign outputDataBuffer_7_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_7_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_7_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_7_data_MPORT_2_addr = outputDataBuffer_7_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_7_data_MPORT_2_data = outputDataBuffer_7_data[outputDataBuffer_7_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_7_data_MPORT_4_data = wr_D_outBuf_7_data;
  assign outputDataBuffer_7_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_7_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_7_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_8_validBit_MPORT_2_addr = outputDataBuffer_8_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_8_validBit_MPORT_2_data =
    outputDataBuffer_8_validBit[outputDataBuffer_8_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_8_validBit_MPORT_4_data = wr_D_outBuf_8_validBit;
  assign outputDataBuffer_8_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_8_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_8_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_8_data_MPORT_2_addr = outputDataBuffer_8_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_8_data_MPORT_2_data = outputDataBuffer_8_data[outputDataBuffer_8_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_8_data_MPORT_4_data = wr_D_outBuf_8_data;
  assign outputDataBuffer_8_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_8_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_8_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_9_validBit_MPORT_2_addr = outputDataBuffer_9_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_9_validBit_MPORT_2_data =
    outputDataBuffer_9_validBit[outputDataBuffer_9_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_9_validBit_MPORT_4_data = wr_D_outBuf_9_validBit;
  assign outputDataBuffer_9_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_9_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_9_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_9_data_MPORT_2_addr = outputDataBuffer_9_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_9_data_MPORT_2_data = outputDataBuffer_9_data[outputDataBuffer_9_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_9_data_MPORT_4_data = wr_D_outBuf_9_data;
  assign outputDataBuffer_9_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_9_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_9_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_10_validBit_MPORT_2_addr = outputDataBuffer_10_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_10_validBit_MPORT_2_data =
    outputDataBuffer_10_validBit[outputDataBuffer_10_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_10_validBit_MPORT_4_data = wr_D_outBuf_10_validBit;
  assign outputDataBuffer_10_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_10_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_10_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_10_data_MPORT_2_addr = outputDataBuffer_10_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_10_data_MPORT_2_data = outputDataBuffer_10_data[outputDataBuffer_10_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_10_data_MPORT_4_data = wr_D_outBuf_10_data;
  assign outputDataBuffer_10_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_10_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_10_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_11_validBit_MPORT_2_addr = outputDataBuffer_11_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_11_validBit_MPORT_2_data =
    outputDataBuffer_11_validBit[outputDataBuffer_11_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_11_validBit_MPORT_4_data = wr_D_outBuf_11_validBit;
  assign outputDataBuffer_11_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_11_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_11_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_11_data_MPORT_2_addr = outputDataBuffer_11_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_11_data_MPORT_2_data = outputDataBuffer_11_data[outputDataBuffer_11_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_11_data_MPORT_4_data = wr_D_outBuf_11_data;
  assign outputDataBuffer_11_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_11_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_11_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_12_validBit_MPORT_2_addr = outputDataBuffer_12_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_12_validBit_MPORT_2_data =
    outputDataBuffer_12_validBit[outputDataBuffer_12_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_12_validBit_MPORT_4_data = wr_D_outBuf_12_validBit;
  assign outputDataBuffer_12_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_12_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_12_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_12_data_MPORT_2_addr = outputDataBuffer_12_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_12_data_MPORT_2_data = outputDataBuffer_12_data[outputDataBuffer_12_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_12_data_MPORT_4_data = wr_D_outBuf_12_data;
  assign outputDataBuffer_12_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_12_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_12_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_13_validBit_MPORT_2_addr = outputDataBuffer_13_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_13_validBit_MPORT_2_data =
    outputDataBuffer_13_validBit[outputDataBuffer_13_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_13_validBit_MPORT_4_data = wr_D_outBuf_13_validBit;
  assign outputDataBuffer_13_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_13_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_13_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_13_data_MPORT_2_addr = outputDataBuffer_13_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_13_data_MPORT_2_data = outputDataBuffer_13_data[outputDataBuffer_13_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_13_data_MPORT_4_data = wr_D_outBuf_13_data;
  assign outputDataBuffer_13_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_13_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_13_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_14_validBit_MPORT_2_addr = outputDataBuffer_14_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_14_validBit_MPORT_2_data =
    outputDataBuffer_14_validBit[outputDataBuffer_14_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_14_validBit_MPORT_4_data = wr_D_outBuf_14_validBit;
  assign outputDataBuffer_14_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_14_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_14_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_14_data_MPORT_2_addr = outputDataBuffer_14_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_14_data_MPORT_2_data = outputDataBuffer_14_data[outputDataBuffer_14_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_14_data_MPORT_4_data = wr_D_outBuf_14_data;
  assign outputDataBuffer_14_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_14_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_14_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_15_validBit_MPORT_2_addr = outputDataBuffer_15_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_15_validBit_MPORT_2_data =
    outputDataBuffer_15_validBit[outputDataBuffer_15_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_15_validBit_MPORT_4_data = wr_D_outBuf_15_validBit;
  assign outputDataBuffer_15_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_15_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_15_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_15_data_MPORT_2_addr = outputDataBuffer_15_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_15_data_MPORT_2_data = outputDataBuffer_15_data[outputDataBuffer_15_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_15_data_MPORT_4_data = wr_D_outBuf_15_data;
  assign outputDataBuffer_15_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_15_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_15_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_16_validBit_MPORT_2_addr = outputDataBuffer_16_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_16_validBit_MPORT_2_data =
    outputDataBuffer_16_validBit[outputDataBuffer_16_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_16_validBit_MPORT_4_data = wr_D_outBuf_16_validBit;
  assign outputDataBuffer_16_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_16_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_16_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_16_data_MPORT_2_addr = outputDataBuffer_16_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_16_data_MPORT_2_data = outputDataBuffer_16_data[outputDataBuffer_16_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_16_data_MPORT_4_data = wr_D_outBuf_16_data;
  assign outputDataBuffer_16_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_16_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_16_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_17_validBit_MPORT_2_addr = outputDataBuffer_17_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_17_validBit_MPORT_2_data =
    outputDataBuffer_17_validBit[outputDataBuffer_17_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_17_validBit_MPORT_4_data = wr_D_outBuf_17_validBit;
  assign outputDataBuffer_17_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_17_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_17_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_17_data_MPORT_2_addr = outputDataBuffer_17_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_17_data_MPORT_2_data = outputDataBuffer_17_data[outputDataBuffer_17_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_17_data_MPORT_4_data = wr_D_outBuf_17_data;
  assign outputDataBuffer_17_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_17_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_17_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_18_validBit_MPORT_2_addr = outputDataBuffer_18_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_18_validBit_MPORT_2_data =
    outputDataBuffer_18_validBit[outputDataBuffer_18_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_18_validBit_MPORT_4_data = wr_D_outBuf_18_validBit;
  assign outputDataBuffer_18_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_18_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_18_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_18_data_MPORT_2_addr = outputDataBuffer_18_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_18_data_MPORT_2_data = outputDataBuffer_18_data[outputDataBuffer_18_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_18_data_MPORT_4_data = wr_D_outBuf_18_data;
  assign outputDataBuffer_18_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_18_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_18_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_19_validBit_MPORT_2_addr = outputDataBuffer_19_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_19_validBit_MPORT_2_data =
    outputDataBuffer_19_validBit[outputDataBuffer_19_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_19_validBit_MPORT_4_data = wr_D_outBuf_19_validBit;
  assign outputDataBuffer_19_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_19_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_19_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_19_data_MPORT_2_addr = outputDataBuffer_19_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_19_data_MPORT_2_data = outputDataBuffer_19_data[outputDataBuffer_19_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_19_data_MPORT_4_data = wr_D_outBuf_19_data;
  assign outputDataBuffer_19_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_19_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_19_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_20_validBit_MPORT_2_addr = outputDataBuffer_20_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_20_validBit_MPORT_2_data =
    outputDataBuffer_20_validBit[outputDataBuffer_20_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_20_validBit_MPORT_4_data = wr_D_outBuf_20_validBit;
  assign outputDataBuffer_20_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_20_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_20_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_20_data_MPORT_2_addr = outputDataBuffer_20_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_20_data_MPORT_2_data = outputDataBuffer_20_data[outputDataBuffer_20_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_20_data_MPORT_4_data = wr_D_outBuf_20_data;
  assign outputDataBuffer_20_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_20_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_20_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_21_validBit_MPORT_2_addr = outputDataBuffer_21_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_21_validBit_MPORT_2_data =
    outputDataBuffer_21_validBit[outputDataBuffer_21_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_21_validBit_MPORT_4_data = wr_D_outBuf_21_validBit;
  assign outputDataBuffer_21_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_21_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_21_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_21_data_MPORT_2_addr = outputDataBuffer_21_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_21_data_MPORT_2_data = outputDataBuffer_21_data[outputDataBuffer_21_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_21_data_MPORT_4_data = wr_D_outBuf_21_data;
  assign outputDataBuffer_21_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_21_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_21_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_22_validBit_MPORT_2_addr = outputDataBuffer_22_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_22_validBit_MPORT_2_data =
    outputDataBuffer_22_validBit[outputDataBuffer_22_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_22_validBit_MPORT_4_data = wr_D_outBuf_22_validBit;
  assign outputDataBuffer_22_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_22_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_22_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_22_data_MPORT_2_addr = outputDataBuffer_22_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_22_data_MPORT_2_data = outputDataBuffer_22_data[outputDataBuffer_22_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_22_data_MPORT_4_data = wr_D_outBuf_22_data;
  assign outputDataBuffer_22_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_22_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_22_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_23_validBit_MPORT_2_addr = outputDataBuffer_23_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_23_validBit_MPORT_2_data =
    outputDataBuffer_23_validBit[outputDataBuffer_23_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_23_validBit_MPORT_4_data = wr_D_outBuf_23_validBit;
  assign outputDataBuffer_23_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_23_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_23_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_23_data_MPORT_2_addr = outputDataBuffer_23_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_23_data_MPORT_2_data = outputDataBuffer_23_data[outputDataBuffer_23_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_23_data_MPORT_4_data = wr_D_outBuf_23_data;
  assign outputDataBuffer_23_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_23_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_23_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_24_validBit_MPORT_2_addr = outputDataBuffer_24_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_24_validBit_MPORT_2_data =
    outputDataBuffer_24_validBit[outputDataBuffer_24_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_24_validBit_MPORT_4_data = wr_D_outBuf_24_validBit;
  assign outputDataBuffer_24_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_24_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_24_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_24_data_MPORT_2_addr = outputDataBuffer_24_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_24_data_MPORT_2_data = outputDataBuffer_24_data[outputDataBuffer_24_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_24_data_MPORT_4_data = wr_D_outBuf_24_data;
  assign outputDataBuffer_24_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_24_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_24_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_25_validBit_MPORT_2_addr = outputDataBuffer_25_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_25_validBit_MPORT_2_data =
    outputDataBuffer_25_validBit[outputDataBuffer_25_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_25_validBit_MPORT_4_data = wr_D_outBuf_25_validBit;
  assign outputDataBuffer_25_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_25_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_25_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_25_data_MPORT_2_addr = outputDataBuffer_25_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_25_data_MPORT_2_data = outputDataBuffer_25_data[outputDataBuffer_25_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_25_data_MPORT_4_data = wr_D_outBuf_25_data;
  assign outputDataBuffer_25_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_25_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_25_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_26_validBit_MPORT_2_addr = outputDataBuffer_26_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_26_validBit_MPORT_2_data =
    outputDataBuffer_26_validBit[outputDataBuffer_26_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_26_validBit_MPORT_4_data = wr_D_outBuf_26_validBit;
  assign outputDataBuffer_26_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_26_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_26_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_26_data_MPORT_2_addr = outputDataBuffer_26_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_26_data_MPORT_2_data = outputDataBuffer_26_data[outputDataBuffer_26_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_26_data_MPORT_4_data = wr_D_outBuf_26_data;
  assign outputDataBuffer_26_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_26_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_26_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_27_validBit_MPORT_2_addr = outputDataBuffer_27_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_27_validBit_MPORT_2_data =
    outputDataBuffer_27_validBit[outputDataBuffer_27_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_27_validBit_MPORT_4_data = wr_D_outBuf_27_validBit;
  assign outputDataBuffer_27_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_27_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_27_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_27_data_MPORT_2_addr = outputDataBuffer_27_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_27_data_MPORT_2_data = outputDataBuffer_27_data[outputDataBuffer_27_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_27_data_MPORT_4_data = wr_D_outBuf_27_data;
  assign outputDataBuffer_27_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_27_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_27_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_28_validBit_MPORT_2_addr = outputDataBuffer_28_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_28_validBit_MPORT_2_data =
    outputDataBuffer_28_validBit[outputDataBuffer_28_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_28_validBit_MPORT_4_data = wr_D_outBuf_28_validBit;
  assign outputDataBuffer_28_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_28_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_28_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_28_data_MPORT_2_addr = outputDataBuffer_28_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_28_data_MPORT_2_data = outputDataBuffer_28_data[outputDataBuffer_28_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_28_data_MPORT_4_data = wr_D_outBuf_28_data;
  assign outputDataBuffer_28_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_28_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_28_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_29_validBit_MPORT_2_addr = outputDataBuffer_29_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_29_validBit_MPORT_2_data =
    outputDataBuffer_29_validBit[outputDataBuffer_29_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_29_validBit_MPORT_4_data = wr_D_outBuf_29_validBit;
  assign outputDataBuffer_29_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_29_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_29_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_29_data_MPORT_2_addr = outputDataBuffer_29_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_29_data_MPORT_2_data = outputDataBuffer_29_data[outputDataBuffer_29_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_29_data_MPORT_4_data = wr_D_outBuf_29_data;
  assign outputDataBuffer_29_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_29_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_29_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_30_validBit_MPORT_2_addr = outputDataBuffer_30_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_30_validBit_MPORT_2_data =
    outputDataBuffer_30_validBit[outputDataBuffer_30_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_30_validBit_MPORT_4_data = wr_D_outBuf_30_validBit;
  assign outputDataBuffer_30_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_30_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_30_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_30_data_MPORT_2_addr = outputDataBuffer_30_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_30_data_MPORT_2_data = outputDataBuffer_30_data[outputDataBuffer_30_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_30_data_MPORT_4_data = wr_D_outBuf_30_data;
  assign outputDataBuffer_30_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_30_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_30_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_31_validBit_MPORT_2_addr = outputDataBuffer_31_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_31_validBit_MPORT_2_data =
    outputDataBuffer_31_validBit[outputDataBuffer_31_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_31_validBit_MPORT_4_data = wr_D_outBuf_31_validBit;
  assign outputDataBuffer_31_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_31_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_31_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_31_data_MPORT_2_addr = outputDataBuffer_31_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_31_data_MPORT_2_data = outputDataBuffer_31_data[outputDataBuffer_31_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_31_data_MPORT_4_data = wr_D_outBuf_31_data;
  assign outputDataBuffer_31_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_31_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_31_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_32_validBit_MPORT_2_addr = outputDataBuffer_32_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_32_validBit_MPORT_2_data =
    outputDataBuffer_32_validBit[outputDataBuffer_32_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_32_validBit_MPORT_4_data = wr_D_outBuf_32_validBit;
  assign outputDataBuffer_32_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_32_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_32_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_32_data_MPORT_2_addr = outputDataBuffer_32_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_32_data_MPORT_2_data = outputDataBuffer_32_data[outputDataBuffer_32_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_32_data_MPORT_4_data = wr_D_outBuf_32_data;
  assign outputDataBuffer_32_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_32_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_32_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_33_validBit_MPORT_2_addr = outputDataBuffer_33_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_33_validBit_MPORT_2_data =
    outputDataBuffer_33_validBit[outputDataBuffer_33_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_33_validBit_MPORT_4_data = wr_D_outBuf_33_validBit;
  assign outputDataBuffer_33_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_33_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_33_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_33_data_MPORT_2_addr = outputDataBuffer_33_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_33_data_MPORT_2_data = outputDataBuffer_33_data[outputDataBuffer_33_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_33_data_MPORT_4_data = wr_D_outBuf_33_data;
  assign outputDataBuffer_33_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_33_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_33_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_34_validBit_MPORT_2_addr = outputDataBuffer_34_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_34_validBit_MPORT_2_data =
    outputDataBuffer_34_validBit[outputDataBuffer_34_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_34_validBit_MPORT_4_data = wr_D_outBuf_34_validBit;
  assign outputDataBuffer_34_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_34_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_34_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_34_data_MPORT_2_addr = outputDataBuffer_34_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_34_data_MPORT_2_data = outputDataBuffer_34_data[outputDataBuffer_34_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_34_data_MPORT_4_data = wr_D_outBuf_34_data;
  assign outputDataBuffer_34_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_34_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_34_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_35_validBit_MPORT_2_addr = outputDataBuffer_35_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_35_validBit_MPORT_2_data =
    outputDataBuffer_35_validBit[outputDataBuffer_35_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_35_validBit_MPORT_4_data = wr_D_outBuf_35_validBit;
  assign outputDataBuffer_35_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_35_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_35_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_35_data_MPORT_2_addr = outputDataBuffer_35_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_35_data_MPORT_2_data = outputDataBuffer_35_data[outputDataBuffer_35_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_35_data_MPORT_4_data = wr_D_outBuf_35_data;
  assign outputDataBuffer_35_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_35_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_35_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_36_validBit_MPORT_2_addr = outputDataBuffer_36_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_36_validBit_MPORT_2_data =
    outputDataBuffer_36_validBit[outputDataBuffer_36_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_36_validBit_MPORT_4_data = wr_D_outBuf_36_validBit;
  assign outputDataBuffer_36_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_36_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_36_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_36_data_MPORT_2_addr = outputDataBuffer_36_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_36_data_MPORT_2_data = outputDataBuffer_36_data[outputDataBuffer_36_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_36_data_MPORT_4_data = wr_D_outBuf_36_data;
  assign outputDataBuffer_36_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_36_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_36_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_37_validBit_MPORT_2_addr = outputDataBuffer_37_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_37_validBit_MPORT_2_data =
    outputDataBuffer_37_validBit[outputDataBuffer_37_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_37_validBit_MPORT_4_data = wr_D_outBuf_37_validBit;
  assign outputDataBuffer_37_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_37_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_37_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_37_data_MPORT_2_addr = outputDataBuffer_37_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_37_data_MPORT_2_data = outputDataBuffer_37_data[outputDataBuffer_37_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_37_data_MPORT_4_data = wr_D_outBuf_37_data;
  assign outputDataBuffer_37_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_37_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_37_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_38_validBit_MPORT_2_addr = outputDataBuffer_38_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_38_validBit_MPORT_2_data =
    outputDataBuffer_38_validBit[outputDataBuffer_38_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_38_validBit_MPORT_4_data = wr_D_outBuf_38_validBit;
  assign outputDataBuffer_38_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_38_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_38_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_38_data_MPORT_2_addr = outputDataBuffer_38_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_38_data_MPORT_2_data = outputDataBuffer_38_data[outputDataBuffer_38_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_38_data_MPORT_4_data = wr_D_outBuf_38_data;
  assign outputDataBuffer_38_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_38_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_38_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_39_validBit_MPORT_2_addr = outputDataBuffer_39_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_39_validBit_MPORT_2_data =
    outputDataBuffer_39_validBit[outputDataBuffer_39_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_39_validBit_MPORT_4_data = wr_D_outBuf_39_validBit;
  assign outputDataBuffer_39_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_39_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_39_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_39_data_MPORT_2_addr = outputDataBuffer_39_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_39_data_MPORT_2_data = outputDataBuffer_39_data[outputDataBuffer_39_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_39_data_MPORT_4_data = wr_D_outBuf_39_data;
  assign outputDataBuffer_39_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_39_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_39_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_40_validBit_MPORT_2_addr = outputDataBuffer_40_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_40_validBit_MPORT_2_data =
    outputDataBuffer_40_validBit[outputDataBuffer_40_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_40_validBit_MPORT_4_data = wr_D_outBuf_40_validBit;
  assign outputDataBuffer_40_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_40_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_40_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_40_data_MPORT_2_addr = outputDataBuffer_40_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_40_data_MPORT_2_data = outputDataBuffer_40_data[outputDataBuffer_40_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_40_data_MPORT_4_data = wr_D_outBuf_40_data;
  assign outputDataBuffer_40_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_40_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_40_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_41_validBit_MPORT_2_addr = outputDataBuffer_41_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_41_validBit_MPORT_2_data =
    outputDataBuffer_41_validBit[outputDataBuffer_41_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_41_validBit_MPORT_4_data = wr_D_outBuf_41_validBit;
  assign outputDataBuffer_41_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_41_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_41_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_41_data_MPORT_2_addr = outputDataBuffer_41_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_41_data_MPORT_2_data = outputDataBuffer_41_data[outputDataBuffer_41_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_41_data_MPORT_4_data = wr_D_outBuf_41_data;
  assign outputDataBuffer_41_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_41_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_41_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_42_validBit_MPORT_2_addr = outputDataBuffer_42_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_42_validBit_MPORT_2_data =
    outputDataBuffer_42_validBit[outputDataBuffer_42_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_42_validBit_MPORT_4_data = wr_D_outBuf_42_validBit;
  assign outputDataBuffer_42_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_42_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_42_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_42_data_MPORT_2_addr = outputDataBuffer_42_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_42_data_MPORT_2_data = outputDataBuffer_42_data[outputDataBuffer_42_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_42_data_MPORT_4_data = wr_D_outBuf_42_data;
  assign outputDataBuffer_42_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_42_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_42_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_43_validBit_MPORT_2_addr = outputDataBuffer_43_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_43_validBit_MPORT_2_data =
    outputDataBuffer_43_validBit[outputDataBuffer_43_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_43_validBit_MPORT_4_data = wr_D_outBuf_43_validBit;
  assign outputDataBuffer_43_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_43_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_43_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_43_data_MPORT_2_addr = outputDataBuffer_43_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_43_data_MPORT_2_data = outputDataBuffer_43_data[outputDataBuffer_43_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_43_data_MPORT_4_data = wr_D_outBuf_43_data;
  assign outputDataBuffer_43_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_43_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_43_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_44_validBit_MPORT_2_addr = outputDataBuffer_44_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_44_validBit_MPORT_2_data =
    outputDataBuffer_44_validBit[outputDataBuffer_44_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_44_validBit_MPORT_4_data = wr_D_outBuf_44_validBit;
  assign outputDataBuffer_44_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_44_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_44_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_44_data_MPORT_2_addr = outputDataBuffer_44_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_44_data_MPORT_2_data = outputDataBuffer_44_data[outputDataBuffer_44_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_44_data_MPORT_4_data = wr_D_outBuf_44_data;
  assign outputDataBuffer_44_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_44_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_44_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_45_validBit_MPORT_2_addr = outputDataBuffer_45_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_45_validBit_MPORT_2_data =
    outputDataBuffer_45_validBit[outputDataBuffer_45_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_45_validBit_MPORT_4_data = wr_D_outBuf_45_validBit;
  assign outputDataBuffer_45_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_45_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_45_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_45_data_MPORT_2_addr = outputDataBuffer_45_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_45_data_MPORT_2_data = outputDataBuffer_45_data[outputDataBuffer_45_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_45_data_MPORT_4_data = wr_D_outBuf_45_data;
  assign outputDataBuffer_45_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_45_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_45_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_46_validBit_MPORT_2_addr = outputDataBuffer_46_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_46_validBit_MPORT_2_data =
    outputDataBuffer_46_validBit[outputDataBuffer_46_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_46_validBit_MPORT_4_data = wr_D_outBuf_46_validBit;
  assign outputDataBuffer_46_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_46_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_46_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_46_data_MPORT_2_addr = outputDataBuffer_46_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_46_data_MPORT_2_data = outputDataBuffer_46_data[outputDataBuffer_46_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_46_data_MPORT_4_data = wr_D_outBuf_46_data;
  assign outputDataBuffer_46_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_46_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_46_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_47_validBit_MPORT_2_addr = outputDataBuffer_47_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_47_validBit_MPORT_2_data =
    outputDataBuffer_47_validBit[outputDataBuffer_47_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_47_validBit_MPORT_4_data = wr_D_outBuf_47_validBit;
  assign outputDataBuffer_47_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_47_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_47_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_47_data_MPORT_2_addr = outputDataBuffer_47_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_47_data_MPORT_2_data = outputDataBuffer_47_data[outputDataBuffer_47_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_47_data_MPORT_4_data = wr_D_outBuf_47_data;
  assign outputDataBuffer_47_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_47_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_47_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_48_validBit_MPORT_2_addr = outputDataBuffer_48_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_48_validBit_MPORT_2_data =
    outputDataBuffer_48_validBit[outputDataBuffer_48_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_48_validBit_MPORT_4_data = wr_D_outBuf_48_validBit;
  assign outputDataBuffer_48_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_48_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_48_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_48_data_MPORT_2_addr = outputDataBuffer_48_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_48_data_MPORT_2_data = outputDataBuffer_48_data[outputDataBuffer_48_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_48_data_MPORT_4_data = wr_D_outBuf_48_data;
  assign outputDataBuffer_48_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_48_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_48_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_49_validBit_MPORT_2_addr = outputDataBuffer_49_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_49_validBit_MPORT_2_data =
    outputDataBuffer_49_validBit[outputDataBuffer_49_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_49_validBit_MPORT_4_data = wr_D_outBuf_49_validBit;
  assign outputDataBuffer_49_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_49_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_49_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_49_data_MPORT_2_addr = outputDataBuffer_49_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_49_data_MPORT_2_data = outputDataBuffer_49_data[outputDataBuffer_49_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_49_data_MPORT_4_data = wr_D_outBuf_49_data;
  assign outputDataBuffer_49_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_49_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_49_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_50_validBit_MPORT_2_addr = outputDataBuffer_50_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_50_validBit_MPORT_2_data =
    outputDataBuffer_50_validBit[outputDataBuffer_50_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_50_validBit_MPORT_4_data = wr_D_outBuf_50_validBit;
  assign outputDataBuffer_50_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_50_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_50_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_50_data_MPORT_2_addr = outputDataBuffer_50_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_50_data_MPORT_2_data = outputDataBuffer_50_data[outputDataBuffer_50_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_50_data_MPORT_4_data = wr_D_outBuf_50_data;
  assign outputDataBuffer_50_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_50_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_50_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_51_validBit_MPORT_2_addr = outputDataBuffer_51_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_51_validBit_MPORT_2_data =
    outputDataBuffer_51_validBit[outputDataBuffer_51_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_51_validBit_MPORT_4_data = wr_D_outBuf_51_validBit;
  assign outputDataBuffer_51_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_51_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_51_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_51_data_MPORT_2_addr = outputDataBuffer_51_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_51_data_MPORT_2_data = outputDataBuffer_51_data[outputDataBuffer_51_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_51_data_MPORT_4_data = wr_D_outBuf_51_data;
  assign outputDataBuffer_51_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_51_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_51_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_52_validBit_MPORT_2_addr = outputDataBuffer_52_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_52_validBit_MPORT_2_data =
    outputDataBuffer_52_validBit[outputDataBuffer_52_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_52_validBit_MPORT_4_data = wr_D_outBuf_52_validBit;
  assign outputDataBuffer_52_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_52_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_52_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_52_data_MPORT_2_addr = outputDataBuffer_52_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_52_data_MPORT_2_data = outputDataBuffer_52_data[outputDataBuffer_52_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_52_data_MPORT_4_data = wr_D_outBuf_52_data;
  assign outputDataBuffer_52_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_52_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_52_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_53_validBit_MPORT_2_addr = outputDataBuffer_53_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_53_validBit_MPORT_2_data =
    outputDataBuffer_53_validBit[outputDataBuffer_53_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_53_validBit_MPORT_4_data = wr_D_outBuf_53_validBit;
  assign outputDataBuffer_53_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_53_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_53_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_53_data_MPORT_2_addr = outputDataBuffer_53_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_53_data_MPORT_2_data = outputDataBuffer_53_data[outputDataBuffer_53_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_53_data_MPORT_4_data = wr_D_outBuf_53_data;
  assign outputDataBuffer_53_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_53_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_53_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_54_validBit_MPORT_2_addr = outputDataBuffer_54_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_54_validBit_MPORT_2_data =
    outputDataBuffer_54_validBit[outputDataBuffer_54_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_54_validBit_MPORT_4_data = wr_D_outBuf_54_validBit;
  assign outputDataBuffer_54_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_54_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_54_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_54_data_MPORT_2_addr = outputDataBuffer_54_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_54_data_MPORT_2_data = outputDataBuffer_54_data[outputDataBuffer_54_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_54_data_MPORT_4_data = wr_D_outBuf_54_data;
  assign outputDataBuffer_54_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_54_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_54_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_55_validBit_MPORT_2_addr = outputDataBuffer_55_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_55_validBit_MPORT_2_data =
    outputDataBuffer_55_validBit[outputDataBuffer_55_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_55_validBit_MPORT_4_data = wr_D_outBuf_55_validBit;
  assign outputDataBuffer_55_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_55_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_55_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_55_data_MPORT_2_addr = outputDataBuffer_55_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_55_data_MPORT_2_data = outputDataBuffer_55_data[outputDataBuffer_55_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_55_data_MPORT_4_data = wr_D_outBuf_55_data;
  assign outputDataBuffer_55_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_55_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_55_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_56_validBit_MPORT_2_addr = outputDataBuffer_56_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_56_validBit_MPORT_2_data =
    outputDataBuffer_56_validBit[outputDataBuffer_56_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_56_validBit_MPORT_4_data = wr_D_outBuf_56_validBit;
  assign outputDataBuffer_56_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_56_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_56_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_56_data_MPORT_2_addr = outputDataBuffer_56_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_56_data_MPORT_2_data = outputDataBuffer_56_data[outputDataBuffer_56_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_56_data_MPORT_4_data = wr_D_outBuf_56_data;
  assign outputDataBuffer_56_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_56_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_56_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_57_validBit_MPORT_2_addr = outputDataBuffer_57_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_57_validBit_MPORT_2_data =
    outputDataBuffer_57_validBit[outputDataBuffer_57_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_57_validBit_MPORT_4_data = wr_D_outBuf_57_validBit;
  assign outputDataBuffer_57_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_57_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_57_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_57_data_MPORT_2_addr = outputDataBuffer_57_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_57_data_MPORT_2_data = outputDataBuffer_57_data[outputDataBuffer_57_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_57_data_MPORT_4_data = wr_D_outBuf_57_data;
  assign outputDataBuffer_57_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_57_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_57_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_58_validBit_MPORT_2_addr = outputDataBuffer_58_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_58_validBit_MPORT_2_data =
    outputDataBuffer_58_validBit[outputDataBuffer_58_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_58_validBit_MPORT_4_data = wr_D_outBuf_58_validBit;
  assign outputDataBuffer_58_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_58_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_58_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_58_data_MPORT_2_addr = outputDataBuffer_58_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_58_data_MPORT_2_data = outputDataBuffer_58_data[outputDataBuffer_58_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_58_data_MPORT_4_data = wr_D_outBuf_58_data;
  assign outputDataBuffer_58_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_58_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_58_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_59_validBit_MPORT_2_addr = outputDataBuffer_59_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_59_validBit_MPORT_2_data =
    outputDataBuffer_59_validBit[outputDataBuffer_59_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_59_validBit_MPORT_4_data = wr_D_outBuf_59_validBit;
  assign outputDataBuffer_59_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_59_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_59_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_59_data_MPORT_2_addr = outputDataBuffer_59_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_59_data_MPORT_2_data = outputDataBuffer_59_data[outputDataBuffer_59_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_59_data_MPORT_4_data = wr_D_outBuf_59_data;
  assign outputDataBuffer_59_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_59_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_59_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_60_validBit_MPORT_2_addr = outputDataBuffer_60_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_60_validBit_MPORT_2_data =
    outputDataBuffer_60_validBit[outputDataBuffer_60_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_60_validBit_MPORT_4_data = wr_D_outBuf_60_validBit;
  assign outputDataBuffer_60_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_60_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_60_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_60_data_MPORT_2_addr = outputDataBuffer_60_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_60_data_MPORT_2_data = outputDataBuffer_60_data[outputDataBuffer_60_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_60_data_MPORT_4_data = wr_D_outBuf_60_data;
  assign outputDataBuffer_60_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_60_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_60_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_61_validBit_MPORT_2_addr = outputDataBuffer_61_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_61_validBit_MPORT_2_data =
    outputDataBuffer_61_validBit[outputDataBuffer_61_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_61_validBit_MPORT_4_data = wr_D_outBuf_61_validBit;
  assign outputDataBuffer_61_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_61_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_61_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_61_data_MPORT_2_addr = outputDataBuffer_61_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_61_data_MPORT_2_data = outputDataBuffer_61_data[outputDataBuffer_61_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_61_data_MPORT_4_data = wr_D_outBuf_61_data;
  assign outputDataBuffer_61_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_61_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_61_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_62_validBit_MPORT_2_addr = outputDataBuffer_62_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_62_validBit_MPORT_2_data =
    outputDataBuffer_62_validBit[outputDataBuffer_62_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_62_validBit_MPORT_4_data = wr_D_outBuf_62_validBit;
  assign outputDataBuffer_62_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_62_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_62_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_62_data_MPORT_2_addr = outputDataBuffer_62_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_62_data_MPORT_2_data = outputDataBuffer_62_data[outputDataBuffer_62_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_62_data_MPORT_4_data = wr_D_outBuf_62_data;
  assign outputDataBuffer_62_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_62_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_62_data_MPORT_4_en = 1'h1;
  assign outputDataBuffer_63_validBit_MPORT_2_addr = outputDataBuffer_63_validBit_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_63_validBit_MPORT_2_data =
    outputDataBuffer_63_validBit[outputDataBuffer_63_validBit_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_63_validBit_MPORT_4_data = wr_D_outBuf_63_validBit;
  assign outputDataBuffer_63_validBit_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_63_validBit_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_63_validBit_MPORT_4_en = 1'h1;
  assign outputDataBuffer_63_data_MPORT_2_addr = outputDataBuffer_63_data_MPORT_2_addr_pipe_0;
  assign outputDataBuffer_63_data_MPORT_2_data = outputDataBuffer_63_data[outputDataBuffer_63_data_MPORT_2_addr]; // @[BP.scala 47:37]
  assign outputDataBuffer_63_data_MPORT_4_data = wr_D_outBuf_63_data;
  assign outputDataBuffer_63_data_MPORT_4_addr = wr_Addr_outBuf;
  assign outputDataBuffer_63_data_MPORT_4_mask = 1'h1;
  assign outputDataBuffer_63_data_MPORT_4_en = 1'h1;
  assign io_rd_D_outBuf_0_validBit = outputDataBuffer_0_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_0_data = outputDataBuffer_0_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_1_validBit = outputDataBuffer_1_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_1_data = outputDataBuffer_1_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_2_validBit = outputDataBuffer_2_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_2_data = outputDataBuffer_2_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_3_validBit = outputDataBuffer_3_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_3_data = outputDataBuffer_3_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_4_validBit = outputDataBuffer_4_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_4_data = outputDataBuffer_4_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_5_validBit = outputDataBuffer_5_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_5_data = outputDataBuffer_5_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_6_validBit = outputDataBuffer_6_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_6_data = outputDataBuffer_6_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_7_validBit = outputDataBuffer_7_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_7_data = outputDataBuffer_7_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_8_validBit = outputDataBuffer_8_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_8_data = outputDataBuffer_8_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_9_validBit = outputDataBuffer_9_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_9_data = outputDataBuffer_9_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_10_validBit = outputDataBuffer_10_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_10_data = outputDataBuffer_10_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_11_validBit = outputDataBuffer_11_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_11_data = outputDataBuffer_11_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_12_validBit = outputDataBuffer_12_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_12_data = outputDataBuffer_12_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_13_validBit = outputDataBuffer_13_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_13_data = outputDataBuffer_13_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_14_validBit = outputDataBuffer_14_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_14_data = outputDataBuffer_14_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_15_validBit = outputDataBuffer_15_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_15_data = outputDataBuffer_15_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_16_validBit = outputDataBuffer_16_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_16_data = outputDataBuffer_16_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_17_validBit = outputDataBuffer_17_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_17_data = outputDataBuffer_17_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_18_validBit = outputDataBuffer_18_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_18_data = outputDataBuffer_18_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_19_validBit = outputDataBuffer_19_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_19_data = outputDataBuffer_19_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_20_validBit = outputDataBuffer_20_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_20_data = outputDataBuffer_20_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_21_validBit = outputDataBuffer_21_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_21_data = outputDataBuffer_21_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_22_validBit = outputDataBuffer_22_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_22_data = outputDataBuffer_22_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_23_validBit = outputDataBuffer_23_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_23_data = outputDataBuffer_23_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_24_validBit = outputDataBuffer_24_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_24_data = outputDataBuffer_24_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_25_validBit = outputDataBuffer_25_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_25_data = outputDataBuffer_25_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_26_validBit = outputDataBuffer_26_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_26_data = outputDataBuffer_26_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_27_validBit = outputDataBuffer_27_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_27_data = outputDataBuffer_27_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_28_validBit = outputDataBuffer_28_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_28_data = outputDataBuffer_28_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_29_validBit = outputDataBuffer_29_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_29_data = outputDataBuffer_29_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_30_validBit = outputDataBuffer_30_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_30_data = outputDataBuffer_30_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_31_validBit = outputDataBuffer_31_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_31_data = outputDataBuffer_31_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_32_validBit = outputDataBuffer_32_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_32_data = outputDataBuffer_32_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_33_validBit = outputDataBuffer_33_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_33_data = outputDataBuffer_33_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_34_validBit = outputDataBuffer_34_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_34_data = outputDataBuffer_34_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_35_validBit = outputDataBuffer_35_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_35_data = outputDataBuffer_35_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_36_validBit = outputDataBuffer_36_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_36_data = outputDataBuffer_36_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_37_validBit = outputDataBuffer_37_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_37_data = outputDataBuffer_37_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_38_validBit = outputDataBuffer_38_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_38_data = outputDataBuffer_38_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_39_validBit = outputDataBuffer_39_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_39_data = outputDataBuffer_39_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_40_validBit = outputDataBuffer_40_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_40_data = outputDataBuffer_40_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_41_validBit = outputDataBuffer_41_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_41_data = outputDataBuffer_41_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_42_validBit = outputDataBuffer_42_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_42_data = outputDataBuffer_42_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_43_validBit = outputDataBuffer_43_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_43_data = outputDataBuffer_43_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_44_validBit = outputDataBuffer_44_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_44_data = outputDataBuffer_44_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_45_validBit = outputDataBuffer_45_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_45_data = outputDataBuffer_45_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_46_validBit = outputDataBuffer_46_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_46_data = outputDataBuffer_46_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_47_validBit = outputDataBuffer_47_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_47_data = outputDataBuffer_47_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_48_validBit = outputDataBuffer_48_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_48_data = outputDataBuffer_48_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_49_validBit = outputDataBuffer_49_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_49_data = outputDataBuffer_49_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_50_validBit = outputDataBuffer_50_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_50_data = outputDataBuffer_50_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_51_validBit = outputDataBuffer_51_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_51_data = outputDataBuffer_51_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_52_validBit = outputDataBuffer_52_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_52_data = outputDataBuffer_52_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_53_validBit = outputDataBuffer_53_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_53_data = outputDataBuffer_53_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_54_validBit = outputDataBuffer_54_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_54_data = outputDataBuffer_54_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_55_validBit = outputDataBuffer_55_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_55_data = outputDataBuffer_55_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_56_validBit = outputDataBuffer_56_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_56_data = outputDataBuffer_56_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_57_validBit = outputDataBuffer_57_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_57_data = outputDataBuffer_57_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_58_validBit = outputDataBuffer_58_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_58_data = outputDataBuffer_58_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_59_validBit = outputDataBuffer_59_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_59_data = outputDataBuffer_59_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_60_validBit = outputDataBuffer_60_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_60_data = outputDataBuffer_60_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_61_validBit = outputDataBuffer_61_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_61_data = outputDataBuffer_61_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_62_validBit = outputDataBuffer_62_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_62_data = outputDataBuffer_62_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_63_validBit = outputDataBuffer_63_validBit_MPORT_2_data; // @[BP.scala 74:18]
  assign io_rd_D_outBuf_63_data = outputDataBuffer_63_data_MPORT_2_data; // @[BP.scala 74:18]
  assign io_PC_out = array_20_io_PC6_out; // @[BP.scala 346:13]
  assign array_0_clock = clock;
  assign array_0_reset = reset;
  assign array_0_io_d_in_0_a = rd_D_inBuf_0_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_0_valid_a = rd_D_inBuf_0_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_0_b = rd_D_inBuf_1_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_0_valid_b = rd_D_inBuf_1_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_1_a = rd_D_inBuf_2_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_1_valid_a = rd_D_inBuf_2_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_1_b = rd_D_inBuf_3_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_1_valid_b = rd_D_inBuf_3_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_2_a = rd_D_inBuf_4_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_2_valid_a = rd_D_inBuf_4_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_2_b = rd_D_inBuf_5_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_2_valid_b = rd_D_inBuf_5_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_3_a = rd_D_inBuf_6_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_3_valid_a = rd_D_inBuf_6_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_3_b = rd_D_inBuf_7_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_3_valid_b = rd_D_inBuf_7_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_4_a = rd_D_inBuf_8_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_4_valid_a = rd_D_inBuf_8_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_4_b = rd_D_inBuf_9_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_4_valid_b = rd_D_inBuf_9_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_5_a = rd_D_inBuf_10_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_5_valid_a = rd_D_inBuf_10_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_5_b = rd_D_inBuf_11_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_5_valid_b = rd_D_inBuf_11_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_6_a = rd_D_inBuf_12_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_6_valid_a = rd_D_inBuf_12_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_6_b = rd_D_inBuf_13_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_6_valid_b = rd_D_inBuf_13_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_7_a = rd_D_inBuf_14_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_7_valid_a = rd_D_inBuf_14_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_7_b = rd_D_inBuf_15_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_7_valid_b = rd_D_inBuf_15_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_8_a = rd_D_inBuf_16_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_8_valid_a = rd_D_inBuf_16_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_8_b = rd_D_inBuf_17_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_8_valid_b = rd_D_inBuf_17_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_9_a = rd_D_inBuf_18_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_9_valid_a = rd_D_inBuf_18_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_9_b = rd_D_inBuf_19_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_9_valid_b = rd_D_inBuf_19_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_10_a = rd_D_inBuf_20_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_10_valid_a = rd_D_inBuf_20_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_10_b = rd_D_inBuf_21_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_10_valid_b = rd_D_inBuf_21_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_11_a = rd_D_inBuf_22_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_11_valid_a = rd_D_inBuf_22_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_11_b = rd_D_inBuf_23_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_11_valid_b = rd_D_inBuf_23_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_12_a = rd_D_inBuf_24_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_12_valid_a = rd_D_inBuf_24_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_12_b = rd_D_inBuf_25_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_12_valid_b = rd_D_inBuf_25_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_13_a = rd_D_inBuf_26_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_13_valid_a = rd_D_inBuf_26_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_13_b = rd_D_inBuf_27_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_13_valid_b = rd_D_inBuf_27_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_14_a = rd_D_inBuf_28_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_14_valid_a = rd_D_inBuf_28_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_14_b = rd_D_inBuf_29_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_14_valid_b = rd_D_inBuf_29_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_15_a = rd_D_inBuf_30_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_15_valid_a = rd_D_inBuf_30_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_15_b = rd_D_inBuf_31_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_15_valid_b = rd_D_inBuf_31_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_16_a = rd_D_inBuf_32_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_16_valid_a = rd_D_inBuf_32_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_16_b = rd_D_inBuf_33_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_16_valid_b = rd_D_inBuf_33_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_17_a = rd_D_inBuf_34_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_17_valid_a = rd_D_inBuf_34_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_17_b = rd_D_inBuf_35_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_17_valid_b = rd_D_inBuf_35_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_18_a = rd_D_inBuf_36_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_18_valid_a = rd_D_inBuf_36_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_18_b = rd_D_inBuf_37_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_18_valid_b = rd_D_inBuf_37_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_19_a = rd_D_inBuf_38_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_19_valid_a = rd_D_inBuf_38_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_19_b = rd_D_inBuf_39_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_19_valid_b = rd_D_inBuf_39_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_20_a = rd_D_inBuf_40_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_20_valid_a = rd_D_inBuf_40_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_20_b = rd_D_inBuf_41_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_20_valid_b = rd_D_inBuf_41_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_21_a = rd_D_inBuf_42_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_21_valid_a = rd_D_inBuf_42_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_21_b = rd_D_inBuf_43_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_21_valid_b = rd_D_inBuf_43_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_22_a = rd_D_inBuf_44_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_22_valid_a = rd_D_inBuf_44_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_22_b = rd_D_inBuf_45_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_22_valid_b = rd_D_inBuf_45_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_23_a = rd_D_inBuf_46_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_23_valid_a = rd_D_inBuf_46_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_23_b = rd_D_inBuf_47_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_23_valid_b = rd_D_inBuf_47_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_24_a = rd_D_inBuf_48_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_24_valid_a = rd_D_inBuf_48_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_24_b = rd_D_inBuf_49_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_24_valid_b = rd_D_inBuf_49_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_25_a = rd_D_inBuf_50_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_25_valid_a = rd_D_inBuf_50_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_25_b = rd_D_inBuf_51_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_25_valid_b = rd_D_inBuf_51_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_26_a = rd_D_inBuf_52_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_26_valid_a = rd_D_inBuf_52_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_26_b = rd_D_inBuf_53_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_26_valid_b = rd_D_inBuf_53_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_27_a = rd_D_inBuf_54_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_27_valid_a = rd_D_inBuf_54_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_27_b = rd_D_inBuf_55_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_27_valid_b = rd_D_inBuf_55_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_28_a = rd_D_inBuf_56_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_28_valid_a = rd_D_inBuf_56_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_28_b = rd_D_inBuf_57_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_28_valid_b = rd_D_inBuf_57_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_29_a = rd_D_inBuf_58_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_29_valid_a = rd_D_inBuf_58_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_29_b = rd_D_inBuf_59_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_29_valid_b = rd_D_inBuf_59_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_30_a = rd_D_inBuf_60_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_30_valid_a = rd_D_inBuf_60_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_30_b = rd_D_inBuf_61_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_30_valid_b = rd_D_inBuf_61_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_d_in_31_a = rd_D_inBuf_62_data; // @[BP.scala 229:18 BP.scala 232:15]
  assign array_0_io_d_in_31_valid_a = rd_D_inBuf_62_validBit; // @[BP.scala 229:18 BP.scala 233:21]
  assign array_0_io_d_in_31_b = rd_D_inBuf_63_data; // @[BP.scala 229:18 BP.scala 234:15]
  assign array_0_io_d_in_31_valid_b = rd_D_inBuf_63_validBit; // @[BP.scala 229:18 BP.scala 235:21]
  assign array_0_io_wr_en_mem1 = io_wr_en_mem1_0; // @[BP.scala 307:26]
  assign array_0_io_wr_en_mem2 = io_wr_en_mem2_0; // @[BP.scala 308:26]
  assign array_0_io_wr_en_mem3 = io_wr_en_mem3_0; // @[BP.scala 309:26]
  assign array_0_io_wr_en_mem4 = io_wr_en_mem4_0; // @[BP.scala 310:26]
  assign array_0_io_wr_en_mem5 = io_wr_en_mem5_0; // @[BP.scala 311:26]
  assign array_0_io_wr_en_mem6 = io_wr_en_mem6_0; // @[BP.scala 312:26]
  assign array_0_io_wr_instr_mem1 = io_wr_instr_mem1_0; // @[BP.scala 313:29]
  assign array_0_io_wr_instr_mem2 = io_wr_instr_mem2_0; // @[BP.scala 314:29]
  assign array_0_io_wr_instr_mem3 = io_wr_instr_mem3_0; // @[BP.scala 315:29]
  assign array_0_io_wr_instr_mem4 = io_wr_instr_mem4_0; // @[BP.scala 316:29]
  assign array_0_io_wr_instr_mem5 = io_wr_instr_mem5_0; // @[BP.scala 317:29]
  assign array_0_io_wr_instr_mem6 = io_wr_instr_mem6_0; // @[BP.scala 318:29]
  assign array_0_io_PC1_in = PCBegin; // @[BP.scala 291:22]
  assign array_0_io_Addr_in = AddrBegin; // @[BP.scala 292:23]
  assign array_1_clock = clock;
  assign array_1_reset = reset;
  assign array_1_io_d_in_0_a = array_0_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_0_valid_a = array_0_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_0_b = array_0_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_0_valid_b = array_0_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_1_a = array_0_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_1_valid_a = array_0_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_1_b = array_0_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_1_valid_b = array_0_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_2_a = array_0_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_2_valid_a = array_0_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_2_b = array_0_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_2_valid_b = array_0_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_3_a = array_0_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_3_valid_a = array_0_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_3_b = array_0_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_3_valid_b = array_0_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_4_a = array_0_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_4_valid_a = array_0_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_4_b = array_0_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_4_valid_b = array_0_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_5_a = array_0_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_5_valid_a = array_0_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_5_b = array_0_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_5_valid_b = array_0_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_6_a = array_0_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_6_valid_a = array_0_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_6_b = array_0_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_6_valid_b = array_0_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_7_a = array_0_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_7_valid_a = array_0_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_7_b = array_0_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_7_valid_b = array_0_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_8_a = array_0_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_8_valid_a = array_0_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_8_b = array_0_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_8_valid_b = array_0_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_9_a = array_0_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_9_valid_a = array_0_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_9_b = array_0_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_9_valid_b = array_0_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_10_a = array_0_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_10_valid_a = array_0_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_10_b = array_0_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_10_valid_b = array_0_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_11_a = array_0_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_11_valid_a = array_0_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_11_b = array_0_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_11_valid_b = array_0_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_12_a = array_0_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_12_valid_a = array_0_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_12_b = array_0_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_12_valid_b = array_0_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_13_a = array_0_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_13_valid_a = array_0_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_13_b = array_0_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_13_valid_b = array_0_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_14_a = array_0_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_14_valid_a = array_0_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_14_b = array_0_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_14_valid_b = array_0_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_15_a = array_0_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_15_valid_a = array_0_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_15_b = array_0_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_15_valid_b = array_0_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_16_a = array_0_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_16_valid_a = array_0_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_16_b = array_0_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_16_valid_b = array_0_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_17_a = array_0_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_17_valid_a = array_0_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_17_b = array_0_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_17_valid_b = array_0_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_18_a = array_0_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_18_valid_a = array_0_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_18_b = array_0_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_18_valid_b = array_0_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_19_a = array_0_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_19_valid_a = array_0_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_19_b = array_0_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_19_valid_b = array_0_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_20_a = array_0_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_20_valid_a = array_0_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_20_b = array_0_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_20_valid_b = array_0_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_21_a = array_0_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_21_valid_a = array_0_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_21_b = array_0_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_21_valid_b = array_0_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_22_a = array_0_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_22_valid_a = array_0_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_22_b = array_0_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_22_valid_b = array_0_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_23_a = array_0_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_23_valid_a = array_0_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_23_b = array_0_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_23_valid_b = array_0_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_24_a = array_0_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_24_valid_a = array_0_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_24_b = array_0_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_24_valid_b = array_0_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_25_a = array_0_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_25_valid_a = array_0_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_25_b = array_0_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_25_valid_b = array_0_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_26_a = array_0_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_26_valid_a = array_0_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_26_b = array_0_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_26_valid_b = array_0_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_27_a = array_0_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_27_valid_a = array_0_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_27_b = array_0_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_27_valid_b = array_0_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_28_a = array_0_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_28_valid_a = array_0_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_28_b = array_0_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_28_valid_b = array_0_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_29_a = array_0_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_29_valid_a = array_0_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_29_b = array_0_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_29_valid_b = array_0_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_30_a = array_0_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_30_valid_a = array_0_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_30_b = array_0_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_30_valid_b = array_0_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_31_a = array_0_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_31_valid_a = array_0_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_1_io_d_in_31_b = array_0_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_1_io_d_in_31_valid_b = array_0_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_1_io_wr_en_mem1 = io_wr_en_mem1_1; // @[BP.scala 325:28]
  assign array_1_io_wr_en_mem2 = io_wr_en_mem2_1; // @[BP.scala 326:28]
  assign array_1_io_wr_en_mem3 = io_wr_en_mem3_1; // @[BP.scala 327:28]
  assign array_1_io_wr_en_mem4 = io_wr_en_mem4_1; // @[BP.scala 328:28]
  assign array_1_io_wr_en_mem5 = io_wr_en_mem5_1; // @[BP.scala 329:28]
  assign array_1_io_wr_en_mem6 = io_wr_en_mem6_1; // @[BP.scala 330:28]
  assign array_1_io_wr_instr_mem1 = io_wr_instr_mem1_1; // @[BP.scala 331:31]
  assign array_1_io_wr_instr_mem2 = io_wr_instr_mem2_1; // @[BP.scala 332:31]
  assign array_1_io_wr_instr_mem3 = io_wr_instr_mem3_1; // @[BP.scala 333:31]
  assign array_1_io_wr_instr_mem4 = io_wr_instr_mem4_1; // @[BP.scala 334:31]
  assign array_1_io_wr_instr_mem5 = io_wr_instr_mem5_1; // @[BP.scala 335:31]
  assign array_1_io_wr_instr_mem6 = io_wr_instr_mem6_1; // @[BP.scala 336:31]
  assign array_1_io_PC1_in = array_0_io_PC6_out; // @[BP.scala 338:24]
  assign array_1_io_Addr_in = array_0_io_Addr_out; // @[BP.scala 339:25]
  assign array_2_clock = clock;
  assign array_2_reset = reset;
  assign array_2_io_d_in_0_a = array_1_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_0_valid_a = array_1_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_0_b = array_1_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_0_valid_b = array_1_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_1_a = array_1_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_1_valid_a = array_1_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_1_b = array_1_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_1_valid_b = array_1_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_2_a = array_1_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_2_valid_a = array_1_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_2_b = array_1_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_2_valid_b = array_1_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_3_a = array_1_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_3_valid_a = array_1_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_3_b = array_1_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_3_valid_b = array_1_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_4_a = array_1_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_4_valid_a = array_1_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_4_b = array_1_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_4_valid_b = array_1_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_5_a = array_1_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_5_valid_a = array_1_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_5_b = array_1_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_5_valid_b = array_1_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_6_a = array_1_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_6_valid_a = array_1_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_6_b = array_1_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_6_valid_b = array_1_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_7_a = array_1_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_7_valid_a = array_1_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_7_b = array_1_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_7_valid_b = array_1_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_8_a = array_1_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_8_valid_a = array_1_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_8_b = array_1_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_8_valid_b = array_1_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_9_a = array_1_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_9_valid_a = array_1_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_9_b = array_1_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_9_valid_b = array_1_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_10_a = array_1_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_10_valid_a = array_1_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_10_b = array_1_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_10_valid_b = array_1_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_11_a = array_1_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_11_valid_a = array_1_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_11_b = array_1_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_11_valid_b = array_1_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_12_a = array_1_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_12_valid_a = array_1_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_12_b = array_1_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_12_valid_b = array_1_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_13_a = array_1_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_13_valid_a = array_1_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_13_b = array_1_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_13_valid_b = array_1_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_14_a = array_1_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_14_valid_a = array_1_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_14_b = array_1_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_14_valid_b = array_1_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_15_a = array_1_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_15_valid_a = array_1_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_15_b = array_1_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_15_valid_b = array_1_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_16_a = array_1_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_16_valid_a = array_1_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_16_b = array_1_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_16_valid_b = array_1_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_17_a = array_1_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_17_valid_a = array_1_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_17_b = array_1_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_17_valid_b = array_1_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_18_a = array_1_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_18_valid_a = array_1_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_18_b = array_1_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_18_valid_b = array_1_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_19_a = array_1_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_19_valid_a = array_1_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_19_b = array_1_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_19_valid_b = array_1_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_20_a = array_1_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_20_valid_a = array_1_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_20_b = array_1_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_20_valid_b = array_1_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_21_a = array_1_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_21_valid_a = array_1_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_21_b = array_1_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_21_valid_b = array_1_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_22_a = array_1_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_22_valid_a = array_1_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_22_b = array_1_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_22_valid_b = array_1_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_23_a = array_1_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_23_valid_a = array_1_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_23_b = array_1_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_23_valid_b = array_1_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_24_a = array_1_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_24_valid_a = array_1_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_24_b = array_1_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_24_valid_b = array_1_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_25_a = array_1_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_25_valid_a = array_1_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_25_b = array_1_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_25_valid_b = array_1_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_26_a = array_1_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_26_valid_a = array_1_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_26_b = array_1_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_26_valid_b = array_1_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_27_a = array_1_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_27_valid_a = array_1_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_27_b = array_1_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_27_valid_b = array_1_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_28_a = array_1_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_28_valid_a = array_1_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_28_b = array_1_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_28_valid_b = array_1_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_29_a = array_1_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_29_valid_a = array_1_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_29_b = array_1_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_29_valid_b = array_1_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_30_a = array_1_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_30_valid_a = array_1_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_30_b = array_1_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_30_valid_b = array_1_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_31_a = array_1_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_31_valid_a = array_1_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_2_io_d_in_31_b = array_1_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_2_io_d_in_31_valid_b = array_1_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_2_io_wr_en_mem1 = io_wr_en_mem1_2; // @[BP.scala 325:28]
  assign array_2_io_wr_en_mem2 = io_wr_en_mem2_2; // @[BP.scala 326:28]
  assign array_2_io_wr_en_mem3 = io_wr_en_mem3_2; // @[BP.scala 327:28]
  assign array_2_io_wr_en_mem4 = io_wr_en_mem4_2; // @[BP.scala 328:28]
  assign array_2_io_wr_en_mem5 = io_wr_en_mem5_2; // @[BP.scala 329:28]
  assign array_2_io_wr_en_mem6 = io_wr_en_mem6_2; // @[BP.scala 330:28]
  assign array_2_io_wr_instr_mem1 = io_wr_instr_mem1_2; // @[BP.scala 331:31]
  assign array_2_io_wr_instr_mem2 = io_wr_instr_mem2_2; // @[BP.scala 332:31]
  assign array_2_io_wr_instr_mem3 = io_wr_instr_mem3_2; // @[BP.scala 333:31]
  assign array_2_io_wr_instr_mem4 = io_wr_instr_mem4_2; // @[BP.scala 334:31]
  assign array_2_io_wr_instr_mem5 = io_wr_instr_mem5_2; // @[BP.scala 335:31]
  assign array_2_io_wr_instr_mem6 = io_wr_instr_mem6_2; // @[BP.scala 336:31]
  assign array_2_io_PC1_in = array_1_io_PC6_out; // @[BP.scala 338:24]
  assign array_2_io_Addr_in = array_1_io_Addr_out; // @[BP.scala 339:25]
  assign array_3_clock = clock;
  assign array_3_reset = reset;
  assign array_3_io_d_in_0_a = array_2_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_0_valid_a = array_2_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_0_b = array_2_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_0_valid_b = array_2_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_1_a = array_2_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_1_valid_a = array_2_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_1_b = array_2_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_1_valid_b = array_2_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_2_a = array_2_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_2_valid_a = array_2_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_2_b = array_2_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_2_valid_b = array_2_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_3_a = array_2_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_3_valid_a = array_2_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_3_b = array_2_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_3_valid_b = array_2_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_4_a = array_2_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_4_valid_a = array_2_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_4_b = array_2_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_4_valid_b = array_2_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_5_a = array_2_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_5_valid_a = array_2_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_5_b = array_2_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_5_valid_b = array_2_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_6_a = array_2_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_6_valid_a = array_2_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_6_b = array_2_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_6_valid_b = array_2_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_7_a = array_2_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_7_valid_a = array_2_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_7_b = array_2_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_7_valid_b = array_2_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_8_a = array_2_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_8_valid_a = array_2_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_8_b = array_2_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_8_valid_b = array_2_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_9_a = array_2_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_9_valid_a = array_2_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_9_b = array_2_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_9_valid_b = array_2_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_10_a = array_2_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_10_valid_a = array_2_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_10_b = array_2_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_10_valid_b = array_2_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_11_a = array_2_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_11_valid_a = array_2_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_11_b = array_2_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_11_valid_b = array_2_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_12_a = array_2_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_12_valid_a = array_2_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_12_b = array_2_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_12_valid_b = array_2_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_13_a = array_2_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_13_valid_a = array_2_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_13_b = array_2_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_13_valid_b = array_2_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_14_a = array_2_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_14_valid_a = array_2_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_14_b = array_2_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_14_valid_b = array_2_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_15_a = array_2_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_15_valid_a = array_2_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_15_b = array_2_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_15_valid_b = array_2_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_16_a = array_2_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_16_valid_a = array_2_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_16_b = array_2_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_16_valid_b = array_2_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_17_a = array_2_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_17_valid_a = array_2_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_17_b = array_2_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_17_valid_b = array_2_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_18_a = array_2_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_18_valid_a = array_2_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_18_b = array_2_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_18_valid_b = array_2_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_19_a = array_2_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_19_valid_a = array_2_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_19_b = array_2_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_19_valid_b = array_2_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_20_a = array_2_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_20_valid_a = array_2_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_20_b = array_2_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_20_valid_b = array_2_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_21_a = array_2_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_21_valid_a = array_2_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_21_b = array_2_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_21_valid_b = array_2_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_22_a = array_2_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_22_valid_a = array_2_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_22_b = array_2_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_22_valid_b = array_2_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_23_a = array_2_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_23_valid_a = array_2_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_23_b = array_2_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_23_valid_b = array_2_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_24_a = array_2_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_24_valid_a = array_2_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_24_b = array_2_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_24_valid_b = array_2_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_25_a = array_2_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_25_valid_a = array_2_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_25_b = array_2_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_25_valid_b = array_2_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_26_a = array_2_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_26_valid_a = array_2_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_26_b = array_2_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_26_valid_b = array_2_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_27_a = array_2_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_27_valid_a = array_2_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_27_b = array_2_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_27_valid_b = array_2_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_28_a = array_2_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_28_valid_a = array_2_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_28_b = array_2_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_28_valid_b = array_2_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_29_a = array_2_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_29_valid_a = array_2_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_29_b = array_2_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_29_valid_b = array_2_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_30_a = array_2_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_30_valid_a = array_2_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_30_b = array_2_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_30_valid_b = array_2_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_31_a = array_2_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_31_valid_a = array_2_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_3_io_d_in_31_b = array_2_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_3_io_d_in_31_valid_b = array_2_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_3_io_wr_en_mem1 = io_wr_en_mem1_3; // @[BP.scala 325:28]
  assign array_3_io_wr_en_mem2 = io_wr_en_mem2_3; // @[BP.scala 326:28]
  assign array_3_io_wr_en_mem3 = io_wr_en_mem3_3; // @[BP.scala 327:28]
  assign array_3_io_wr_en_mem4 = io_wr_en_mem4_3; // @[BP.scala 328:28]
  assign array_3_io_wr_en_mem5 = io_wr_en_mem5_3; // @[BP.scala 329:28]
  assign array_3_io_wr_en_mem6 = io_wr_en_mem6_3; // @[BP.scala 330:28]
  assign array_3_io_wr_instr_mem1 = io_wr_instr_mem1_3; // @[BP.scala 331:31]
  assign array_3_io_wr_instr_mem2 = io_wr_instr_mem2_3; // @[BP.scala 332:31]
  assign array_3_io_wr_instr_mem3 = io_wr_instr_mem3_3; // @[BP.scala 333:31]
  assign array_3_io_wr_instr_mem4 = io_wr_instr_mem4_3; // @[BP.scala 334:31]
  assign array_3_io_wr_instr_mem5 = io_wr_instr_mem5_3; // @[BP.scala 335:31]
  assign array_3_io_wr_instr_mem6 = io_wr_instr_mem6_3; // @[BP.scala 336:31]
  assign array_3_io_PC1_in = array_2_io_PC6_out; // @[BP.scala 338:24]
  assign array_3_io_Addr_in = array_2_io_Addr_out; // @[BP.scala 339:25]
  assign array_4_clock = clock;
  assign array_4_reset = reset;
  assign array_4_io_d_in_0_a = array_3_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_0_valid_a = array_3_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_0_b = array_3_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_0_valid_b = array_3_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_1_a = array_3_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_1_valid_a = array_3_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_1_b = array_3_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_1_valid_b = array_3_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_2_a = array_3_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_2_valid_a = array_3_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_2_b = array_3_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_2_valid_b = array_3_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_3_a = array_3_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_3_valid_a = array_3_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_3_b = array_3_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_3_valid_b = array_3_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_4_a = array_3_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_4_valid_a = array_3_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_4_b = array_3_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_4_valid_b = array_3_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_5_a = array_3_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_5_valid_a = array_3_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_5_b = array_3_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_5_valid_b = array_3_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_6_a = array_3_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_6_valid_a = array_3_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_6_b = array_3_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_6_valid_b = array_3_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_7_a = array_3_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_7_valid_a = array_3_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_7_b = array_3_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_7_valid_b = array_3_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_8_a = array_3_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_8_valid_a = array_3_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_8_b = array_3_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_8_valid_b = array_3_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_9_a = array_3_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_9_valid_a = array_3_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_9_b = array_3_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_9_valid_b = array_3_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_10_a = array_3_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_10_valid_a = array_3_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_10_b = array_3_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_10_valid_b = array_3_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_11_a = array_3_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_11_valid_a = array_3_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_11_b = array_3_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_11_valid_b = array_3_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_12_a = array_3_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_12_valid_a = array_3_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_12_b = array_3_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_12_valid_b = array_3_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_13_a = array_3_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_13_valid_a = array_3_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_13_b = array_3_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_13_valid_b = array_3_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_14_a = array_3_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_14_valid_a = array_3_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_14_b = array_3_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_14_valid_b = array_3_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_15_a = array_3_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_15_valid_a = array_3_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_15_b = array_3_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_15_valid_b = array_3_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_16_a = array_3_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_16_valid_a = array_3_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_16_b = array_3_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_16_valid_b = array_3_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_17_a = array_3_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_17_valid_a = array_3_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_17_b = array_3_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_17_valid_b = array_3_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_18_a = array_3_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_18_valid_a = array_3_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_18_b = array_3_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_18_valid_b = array_3_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_19_a = array_3_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_19_valid_a = array_3_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_19_b = array_3_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_19_valid_b = array_3_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_20_a = array_3_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_20_valid_a = array_3_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_20_b = array_3_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_20_valid_b = array_3_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_21_a = array_3_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_21_valid_a = array_3_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_21_b = array_3_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_21_valid_b = array_3_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_22_a = array_3_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_22_valid_a = array_3_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_22_b = array_3_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_22_valid_b = array_3_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_23_a = array_3_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_23_valid_a = array_3_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_23_b = array_3_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_23_valid_b = array_3_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_24_a = array_3_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_24_valid_a = array_3_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_24_b = array_3_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_24_valid_b = array_3_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_25_a = array_3_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_25_valid_a = array_3_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_25_b = array_3_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_25_valid_b = array_3_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_26_a = array_3_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_26_valid_a = array_3_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_26_b = array_3_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_26_valid_b = array_3_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_27_a = array_3_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_27_valid_a = array_3_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_27_b = array_3_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_27_valid_b = array_3_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_28_a = array_3_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_28_valid_a = array_3_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_28_b = array_3_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_28_valid_b = array_3_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_29_a = array_3_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_29_valid_a = array_3_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_29_b = array_3_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_29_valid_b = array_3_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_30_a = array_3_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_30_valid_a = array_3_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_30_b = array_3_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_30_valid_b = array_3_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_31_a = array_3_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_31_valid_a = array_3_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_4_io_d_in_31_b = array_3_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_4_io_d_in_31_valid_b = array_3_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_4_io_wr_en_mem1 = io_wr_en_mem1_4; // @[BP.scala 325:28]
  assign array_4_io_wr_en_mem2 = io_wr_en_mem2_4; // @[BP.scala 326:28]
  assign array_4_io_wr_en_mem3 = io_wr_en_mem3_4; // @[BP.scala 327:28]
  assign array_4_io_wr_en_mem4 = io_wr_en_mem4_4; // @[BP.scala 328:28]
  assign array_4_io_wr_en_mem5 = io_wr_en_mem5_4; // @[BP.scala 329:28]
  assign array_4_io_wr_en_mem6 = io_wr_en_mem6_4; // @[BP.scala 330:28]
  assign array_4_io_wr_instr_mem1 = io_wr_instr_mem1_4; // @[BP.scala 331:31]
  assign array_4_io_wr_instr_mem2 = io_wr_instr_mem2_4; // @[BP.scala 332:31]
  assign array_4_io_wr_instr_mem3 = io_wr_instr_mem3_4; // @[BP.scala 333:31]
  assign array_4_io_wr_instr_mem4 = io_wr_instr_mem4_4; // @[BP.scala 334:31]
  assign array_4_io_wr_instr_mem5 = io_wr_instr_mem5_4; // @[BP.scala 335:31]
  assign array_4_io_wr_instr_mem6 = io_wr_instr_mem6_4; // @[BP.scala 336:31]
  assign array_4_io_PC1_in = array_3_io_PC6_out; // @[BP.scala 338:24]
  assign array_4_io_Addr_in = array_3_io_Addr_out; // @[BP.scala 339:25]
  assign array_5_clock = clock;
  assign array_5_reset = reset;
  assign array_5_io_d_in_0_a = array_4_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_0_valid_a = array_4_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_0_b = array_4_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_0_valid_b = array_4_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_1_a = array_4_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_1_valid_a = array_4_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_1_b = array_4_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_1_valid_b = array_4_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_2_a = array_4_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_2_valid_a = array_4_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_2_b = array_4_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_2_valid_b = array_4_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_3_a = array_4_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_3_valid_a = array_4_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_3_b = array_4_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_3_valid_b = array_4_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_4_a = array_4_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_4_valid_a = array_4_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_4_b = array_4_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_4_valid_b = array_4_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_5_a = array_4_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_5_valid_a = array_4_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_5_b = array_4_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_5_valid_b = array_4_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_6_a = array_4_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_6_valid_a = array_4_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_6_b = array_4_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_6_valid_b = array_4_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_7_a = array_4_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_7_valid_a = array_4_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_7_b = array_4_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_7_valid_b = array_4_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_8_a = array_4_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_8_valid_a = array_4_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_8_b = array_4_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_8_valid_b = array_4_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_9_a = array_4_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_9_valid_a = array_4_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_9_b = array_4_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_9_valid_b = array_4_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_10_a = array_4_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_10_valid_a = array_4_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_10_b = array_4_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_10_valid_b = array_4_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_11_a = array_4_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_11_valid_a = array_4_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_11_b = array_4_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_11_valid_b = array_4_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_12_a = array_4_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_12_valid_a = array_4_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_12_b = array_4_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_12_valid_b = array_4_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_13_a = array_4_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_13_valid_a = array_4_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_13_b = array_4_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_13_valid_b = array_4_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_14_a = array_4_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_14_valid_a = array_4_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_14_b = array_4_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_14_valid_b = array_4_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_15_a = array_4_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_15_valid_a = array_4_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_15_b = array_4_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_15_valid_b = array_4_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_16_a = array_4_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_16_valid_a = array_4_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_16_b = array_4_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_16_valid_b = array_4_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_17_a = array_4_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_17_valid_a = array_4_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_17_b = array_4_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_17_valid_b = array_4_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_18_a = array_4_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_18_valid_a = array_4_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_18_b = array_4_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_18_valid_b = array_4_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_19_a = array_4_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_19_valid_a = array_4_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_19_b = array_4_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_19_valid_b = array_4_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_20_a = array_4_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_20_valid_a = array_4_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_20_b = array_4_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_20_valid_b = array_4_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_21_a = array_4_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_21_valid_a = array_4_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_21_b = array_4_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_21_valid_b = array_4_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_22_a = array_4_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_22_valid_a = array_4_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_22_b = array_4_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_22_valid_b = array_4_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_23_a = array_4_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_23_valid_a = array_4_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_23_b = array_4_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_23_valid_b = array_4_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_24_a = array_4_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_24_valid_a = array_4_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_24_b = array_4_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_24_valid_b = array_4_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_25_a = array_4_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_25_valid_a = array_4_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_25_b = array_4_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_25_valid_b = array_4_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_26_a = array_4_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_26_valid_a = array_4_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_26_b = array_4_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_26_valid_b = array_4_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_27_a = array_4_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_27_valid_a = array_4_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_27_b = array_4_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_27_valid_b = array_4_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_28_a = array_4_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_28_valid_a = array_4_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_28_b = array_4_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_28_valid_b = array_4_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_29_a = array_4_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_29_valid_a = array_4_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_29_b = array_4_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_29_valid_b = array_4_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_30_a = array_4_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_30_valid_a = array_4_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_30_b = array_4_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_30_valid_b = array_4_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_31_a = array_4_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_31_valid_a = array_4_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_5_io_d_in_31_b = array_4_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_5_io_d_in_31_valid_b = array_4_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_5_io_wr_en_mem1 = io_wr_en_mem1_5; // @[BP.scala 325:28]
  assign array_5_io_wr_en_mem2 = io_wr_en_mem2_5; // @[BP.scala 326:28]
  assign array_5_io_wr_en_mem3 = io_wr_en_mem3_5; // @[BP.scala 327:28]
  assign array_5_io_wr_en_mem4 = io_wr_en_mem4_5; // @[BP.scala 328:28]
  assign array_5_io_wr_en_mem5 = io_wr_en_mem5_5; // @[BP.scala 329:28]
  assign array_5_io_wr_en_mem6 = io_wr_en_mem6_5; // @[BP.scala 330:28]
  assign array_5_io_wr_instr_mem1 = io_wr_instr_mem1_5; // @[BP.scala 331:31]
  assign array_5_io_wr_instr_mem2 = io_wr_instr_mem2_5; // @[BP.scala 332:31]
  assign array_5_io_wr_instr_mem3 = io_wr_instr_mem3_5; // @[BP.scala 333:31]
  assign array_5_io_wr_instr_mem4 = io_wr_instr_mem4_5; // @[BP.scala 334:31]
  assign array_5_io_wr_instr_mem5 = io_wr_instr_mem5_5; // @[BP.scala 335:31]
  assign array_5_io_wr_instr_mem6 = io_wr_instr_mem6_5; // @[BP.scala 336:31]
  assign array_5_io_PC1_in = array_4_io_PC6_out; // @[BP.scala 338:24]
  assign array_5_io_Addr_in = array_4_io_Addr_out; // @[BP.scala 339:25]
  assign array_6_clock = clock;
  assign array_6_reset = reset;
  assign array_6_io_d_in_0_a = array_5_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_0_valid_a = array_5_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_0_b = array_5_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_0_valid_b = array_5_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_1_a = array_5_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_1_valid_a = array_5_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_1_b = array_5_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_1_valid_b = array_5_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_2_a = array_5_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_2_valid_a = array_5_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_2_b = array_5_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_2_valid_b = array_5_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_3_a = array_5_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_3_valid_a = array_5_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_3_b = array_5_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_3_valid_b = array_5_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_4_a = array_5_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_4_valid_a = array_5_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_4_b = array_5_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_4_valid_b = array_5_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_5_a = array_5_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_5_valid_a = array_5_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_5_b = array_5_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_5_valid_b = array_5_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_6_a = array_5_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_6_valid_a = array_5_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_6_b = array_5_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_6_valid_b = array_5_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_7_a = array_5_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_7_valid_a = array_5_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_7_b = array_5_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_7_valid_b = array_5_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_8_a = array_5_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_8_valid_a = array_5_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_8_b = array_5_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_8_valid_b = array_5_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_9_a = array_5_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_9_valid_a = array_5_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_9_b = array_5_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_9_valid_b = array_5_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_10_a = array_5_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_10_valid_a = array_5_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_10_b = array_5_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_10_valid_b = array_5_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_11_a = array_5_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_11_valid_a = array_5_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_11_b = array_5_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_11_valid_b = array_5_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_12_a = array_5_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_12_valid_a = array_5_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_12_b = array_5_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_12_valid_b = array_5_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_13_a = array_5_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_13_valid_a = array_5_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_13_b = array_5_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_13_valid_b = array_5_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_14_a = array_5_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_14_valid_a = array_5_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_14_b = array_5_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_14_valid_b = array_5_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_15_a = array_5_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_15_valid_a = array_5_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_15_b = array_5_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_15_valid_b = array_5_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_16_a = array_5_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_16_valid_a = array_5_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_16_b = array_5_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_16_valid_b = array_5_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_17_a = array_5_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_17_valid_a = array_5_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_17_b = array_5_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_17_valid_b = array_5_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_18_a = array_5_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_18_valid_a = array_5_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_18_b = array_5_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_18_valid_b = array_5_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_19_a = array_5_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_19_valid_a = array_5_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_19_b = array_5_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_19_valid_b = array_5_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_20_a = array_5_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_20_valid_a = array_5_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_20_b = array_5_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_20_valid_b = array_5_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_21_a = array_5_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_21_valid_a = array_5_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_21_b = array_5_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_21_valid_b = array_5_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_22_a = array_5_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_22_valid_a = array_5_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_22_b = array_5_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_22_valid_b = array_5_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_23_a = array_5_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_23_valid_a = array_5_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_23_b = array_5_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_23_valid_b = array_5_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_24_a = array_5_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_24_valid_a = array_5_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_24_b = array_5_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_24_valid_b = array_5_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_25_a = array_5_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_25_valid_a = array_5_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_25_b = array_5_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_25_valid_b = array_5_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_26_a = array_5_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_26_valid_a = array_5_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_26_b = array_5_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_26_valid_b = array_5_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_27_a = array_5_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_27_valid_a = array_5_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_27_b = array_5_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_27_valid_b = array_5_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_28_a = array_5_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_28_valid_a = array_5_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_28_b = array_5_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_28_valid_b = array_5_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_29_a = array_5_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_29_valid_a = array_5_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_29_b = array_5_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_29_valid_b = array_5_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_30_a = array_5_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_30_valid_a = array_5_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_30_b = array_5_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_30_valid_b = array_5_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_31_a = array_5_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_31_valid_a = array_5_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_6_io_d_in_31_b = array_5_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_6_io_d_in_31_valid_b = array_5_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_6_io_wr_en_mem1 = io_wr_en_mem1_6; // @[BP.scala 325:28]
  assign array_6_io_wr_en_mem2 = io_wr_en_mem2_6; // @[BP.scala 326:28]
  assign array_6_io_wr_en_mem3 = io_wr_en_mem3_6; // @[BP.scala 327:28]
  assign array_6_io_wr_en_mem4 = io_wr_en_mem4_6; // @[BP.scala 328:28]
  assign array_6_io_wr_en_mem5 = io_wr_en_mem5_6; // @[BP.scala 329:28]
  assign array_6_io_wr_en_mem6 = io_wr_en_mem6_6; // @[BP.scala 330:28]
  assign array_6_io_wr_instr_mem1 = io_wr_instr_mem1_6; // @[BP.scala 331:31]
  assign array_6_io_wr_instr_mem2 = io_wr_instr_mem2_6; // @[BP.scala 332:31]
  assign array_6_io_wr_instr_mem3 = io_wr_instr_mem3_6; // @[BP.scala 333:31]
  assign array_6_io_wr_instr_mem4 = io_wr_instr_mem4_6; // @[BP.scala 334:31]
  assign array_6_io_wr_instr_mem5 = io_wr_instr_mem5_6; // @[BP.scala 335:31]
  assign array_6_io_wr_instr_mem6 = io_wr_instr_mem6_6; // @[BP.scala 336:31]
  assign array_6_io_PC1_in = array_5_io_PC6_out; // @[BP.scala 338:24]
  assign array_6_io_Addr_in = array_5_io_Addr_out; // @[BP.scala 339:25]
  assign array_7_clock = clock;
  assign array_7_reset = reset;
  assign array_7_io_d_in_0_a = array_6_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_0_valid_a = array_6_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_0_b = array_6_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_0_valid_b = array_6_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_1_a = array_6_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_1_valid_a = array_6_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_1_b = array_6_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_1_valid_b = array_6_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_2_a = array_6_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_2_valid_a = array_6_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_2_b = array_6_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_2_valid_b = array_6_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_3_a = array_6_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_3_valid_a = array_6_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_3_b = array_6_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_3_valid_b = array_6_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_4_a = array_6_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_4_valid_a = array_6_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_4_b = array_6_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_4_valid_b = array_6_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_5_a = array_6_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_5_valid_a = array_6_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_5_b = array_6_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_5_valid_b = array_6_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_6_a = array_6_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_6_valid_a = array_6_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_6_b = array_6_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_6_valid_b = array_6_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_7_a = array_6_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_7_valid_a = array_6_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_7_b = array_6_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_7_valid_b = array_6_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_8_a = array_6_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_8_valid_a = array_6_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_8_b = array_6_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_8_valid_b = array_6_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_9_a = array_6_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_9_valid_a = array_6_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_9_b = array_6_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_9_valid_b = array_6_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_10_a = array_6_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_10_valid_a = array_6_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_10_b = array_6_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_10_valid_b = array_6_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_11_a = array_6_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_11_valid_a = array_6_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_11_b = array_6_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_11_valid_b = array_6_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_12_a = array_6_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_12_valid_a = array_6_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_12_b = array_6_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_12_valid_b = array_6_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_13_a = array_6_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_13_valid_a = array_6_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_13_b = array_6_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_13_valid_b = array_6_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_14_a = array_6_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_14_valid_a = array_6_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_14_b = array_6_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_14_valid_b = array_6_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_15_a = array_6_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_15_valid_a = array_6_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_15_b = array_6_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_15_valid_b = array_6_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_16_a = array_6_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_16_valid_a = array_6_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_16_b = array_6_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_16_valid_b = array_6_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_17_a = array_6_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_17_valid_a = array_6_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_17_b = array_6_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_17_valid_b = array_6_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_18_a = array_6_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_18_valid_a = array_6_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_18_b = array_6_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_18_valid_b = array_6_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_19_a = array_6_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_19_valid_a = array_6_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_19_b = array_6_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_19_valid_b = array_6_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_20_a = array_6_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_20_valid_a = array_6_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_20_b = array_6_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_20_valid_b = array_6_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_21_a = array_6_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_21_valid_a = array_6_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_21_b = array_6_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_21_valid_b = array_6_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_22_a = array_6_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_22_valid_a = array_6_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_22_b = array_6_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_22_valid_b = array_6_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_23_a = array_6_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_23_valid_a = array_6_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_23_b = array_6_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_23_valid_b = array_6_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_24_a = array_6_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_24_valid_a = array_6_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_24_b = array_6_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_24_valid_b = array_6_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_25_a = array_6_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_25_valid_a = array_6_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_25_b = array_6_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_25_valid_b = array_6_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_26_a = array_6_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_26_valid_a = array_6_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_26_b = array_6_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_26_valid_b = array_6_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_27_a = array_6_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_27_valid_a = array_6_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_27_b = array_6_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_27_valid_b = array_6_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_28_a = array_6_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_28_valid_a = array_6_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_28_b = array_6_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_28_valid_b = array_6_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_29_a = array_6_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_29_valid_a = array_6_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_29_b = array_6_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_29_valid_b = array_6_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_30_a = array_6_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_30_valid_a = array_6_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_30_b = array_6_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_30_valid_b = array_6_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_31_a = array_6_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_31_valid_a = array_6_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_7_io_d_in_31_b = array_6_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_7_io_d_in_31_valid_b = array_6_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_7_io_wr_en_mem1 = io_wr_en_mem1_7; // @[BP.scala 325:28]
  assign array_7_io_wr_en_mem2 = io_wr_en_mem2_7; // @[BP.scala 326:28]
  assign array_7_io_wr_en_mem3 = io_wr_en_mem3_7; // @[BP.scala 327:28]
  assign array_7_io_wr_en_mem4 = io_wr_en_mem4_7; // @[BP.scala 328:28]
  assign array_7_io_wr_en_mem5 = io_wr_en_mem5_7; // @[BP.scala 329:28]
  assign array_7_io_wr_en_mem6 = io_wr_en_mem6_7; // @[BP.scala 330:28]
  assign array_7_io_wr_instr_mem1 = io_wr_instr_mem1_7; // @[BP.scala 331:31]
  assign array_7_io_wr_instr_mem2 = io_wr_instr_mem2_7; // @[BP.scala 332:31]
  assign array_7_io_wr_instr_mem3 = io_wr_instr_mem3_7; // @[BP.scala 333:31]
  assign array_7_io_wr_instr_mem4 = io_wr_instr_mem4_7; // @[BP.scala 334:31]
  assign array_7_io_wr_instr_mem5 = io_wr_instr_mem5_7; // @[BP.scala 335:31]
  assign array_7_io_wr_instr_mem6 = io_wr_instr_mem6_7; // @[BP.scala 336:31]
  assign array_7_io_PC1_in = array_6_io_PC6_out; // @[BP.scala 338:24]
  assign array_7_io_Addr_in = array_6_io_Addr_out; // @[BP.scala 339:25]
  assign array_8_clock = clock;
  assign array_8_reset = reset;
  assign array_8_io_d_in_0_a = array_7_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_0_valid_a = array_7_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_0_b = array_7_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_0_valid_b = array_7_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_1_a = array_7_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_1_valid_a = array_7_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_1_b = array_7_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_1_valid_b = array_7_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_2_a = array_7_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_2_valid_a = array_7_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_2_b = array_7_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_2_valid_b = array_7_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_3_a = array_7_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_3_valid_a = array_7_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_3_b = array_7_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_3_valid_b = array_7_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_4_a = array_7_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_4_valid_a = array_7_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_4_b = array_7_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_4_valid_b = array_7_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_5_a = array_7_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_5_valid_a = array_7_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_5_b = array_7_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_5_valid_b = array_7_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_6_a = array_7_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_6_valid_a = array_7_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_6_b = array_7_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_6_valid_b = array_7_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_7_a = array_7_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_7_valid_a = array_7_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_7_b = array_7_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_7_valid_b = array_7_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_8_a = array_7_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_8_valid_a = array_7_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_8_b = array_7_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_8_valid_b = array_7_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_9_a = array_7_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_9_valid_a = array_7_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_9_b = array_7_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_9_valid_b = array_7_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_10_a = array_7_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_10_valid_a = array_7_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_10_b = array_7_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_10_valid_b = array_7_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_11_a = array_7_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_11_valid_a = array_7_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_11_b = array_7_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_11_valid_b = array_7_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_12_a = array_7_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_12_valid_a = array_7_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_12_b = array_7_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_12_valid_b = array_7_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_13_a = array_7_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_13_valid_a = array_7_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_13_b = array_7_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_13_valid_b = array_7_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_14_a = array_7_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_14_valid_a = array_7_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_14_b = array_7_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_14_valid_b = array_7_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_15_a = array_7_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_15_valid_a = array_7_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_15_b = array_7_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_15_valid_b = array_7_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_16_a = array_7_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_16_valid_a = array_7_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_16_b = array_7_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_16_valid_b = array_7_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_17_a = array_7_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_17_valid_a = array_7_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_17_b = array_7_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_17_valid_b = array_7_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_18_a = array_7_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_18_valid_a = array_7_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_18_b = array_7_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_18_valid_b = array_7_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_19_a = array_7_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_19_valid_a = array_7_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_19_b = array_7_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_19_valid_b = array_7_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_20_a = array_7_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_20_valid_a = array_7_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_20_b = array_7_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_20_valid_b = array_7_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_21_a = array_7_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_21_valid_a = array_7_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_21_b = array_7_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_21_valid_b = array_7_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_22_a = array_7_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_22_valid_a = array_7_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_22_b = array_7_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_22_valid_b = array_7_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_23_a = array_7_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_23_valid_a = array_7_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_23_b = array_7_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_23_valid_b = array_7_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_24_a = array_7_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_24_valid_a = array_7_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_24_b = array_7_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_24_valid_b = array_7_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_25_a = array_7_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_25_valid_a = array_7_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_25_b = array_7_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_25_valid_b = array_7_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_26_a = array_7_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_26_valid_a = array_7_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_26_b = array_7_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_26_valid_b = array_7_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_27_a = array_7_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_27_valid_a = array_7_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_27_b = array_7_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_27_valid_b = array_7_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_28_a = array_7_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_28_valid_a = array_7_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_28_b = array_7_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_28_valid_b = array_7_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_29_a = array_7_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_29_valid_a = array_7_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_29_b = array_7_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_29_valid_b = array_7_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_30_a = array_7_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_30_valid_a = array_7_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_30_b = array_7_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_30_valid_b = array_7_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_31_a = array_7_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_31_valid_a = array_7_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_8_io_d_in_31_b = array_7_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_8_io_d_in_31_valid_b = array_7_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_8_io_wr_en_mem1 = io_wr_en_mem1_8; // @[BP.scala 325:28]
  assign array_8_io_wr_en_mem2 = io_wr_en_mem2_8; // @[BP.scala 326:28]
  assign array_8_io_wr_en_mem3 = io_wr_en_mem3_8; // @[BP.scala 327:28]
  assign array_8_io_wr_en_mem4 = io_wr_en_mem4_8; // @[BP.scala 328:28]
  assign array_8_io_wr_en_mem5 = io_wr_en_mem5_8; // @[BP.scala 329:28]
  assign array_8_io_wr_en_mem6 = io_wr_en_mem6_8; // @[BP.scala 330:28]
  assign array_8_io_wr_instr_mem1 = io_wr_instr_mem1_8; // @[BP.scala 331:31]
  assign array_8_io_wr_instr_mem2 = io_wr_instr_mem2_8; // @[BP.scala 332:31]
  assign array_8_io_wr_instr_mem3 = io_wr_instr_mem3_8; // @[BP.scala 333:31]
  assign array_8_io_wr_instr_mem4 = io_wr_instr_mem4_8; // @[BP.scala 334:31]
  assign array_8_io_wr_instr_mem5 = io_wr_instr_mem5_8; // @[BP.scala 335:31]
  assign array_8_io_wr_instr_mem6 = io_wr_instr_mem6_8; // @[BP.scala 336:31]
  assign array_8_io_PC1_in = array_7_io_PC6_out; // @[BP.scala 338:24]
  assign array_8_io_Addr_in = array_7_io_Addr_out; // @[BP.scala 339:25]
  assign array_9_clock = clock;
  assign array_9_reset = reset;
  assign array_9_io_d_in_0_a = array_8_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_0_valid_a = array_8_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_0_b = array_8_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_0_valid_b = array_8_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_1_a = array_8_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_1_valid_a = array_8_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_1_b = array_8_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_1_valid_b = array_8_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_2_a = array_8_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_2_valid_a = array_8_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_2_b = array_8_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_2_valid_b = array_8_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_3_a = array_8_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_3_valid_a = array_8_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_3_b = array_8_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_3_valid_b = array_8_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_4_a = array_8_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_4_valid_a = array_8_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_4_b = array_8_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_4_valid_b = array_8_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_5_a = array_8_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_5_valid_a = array_8_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_5_b = array_8_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_5_valid_b = array_8_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_6_a = array_8_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_6_valid_a = array_8_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_6_b = array_8_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_6_valid_b = array_8_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_7_a = array_8_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_7_valid_a = array_8_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_7_b = array_8_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_7_valid_b = array_8_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_8_a = array_8_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_8_valid_a = array_8_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_8_b = array_8_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_8_valid_b = array_8_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_9_a = array_8_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_9_valid_a = array_8_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_9_b = array_8_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_9_valid_b = array_8_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_10_a = array_8_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_10_valid_a = array_8_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_10_b = array_8_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_10_valid_b = array_8_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_11_a = array_8_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_11_valid_a = array_8_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_11_b = array_8_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_11_valid_b = array_8_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_12_a = array_8_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_12_valid_a = array_8_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_12_b = array_8_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_12_valid_b = array_8_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_13_a = array_8_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_13_valid_a = array_8_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_13_b = array_8_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_13_valid_b = array_8_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_14_a = array_8_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_14_valid_a = array_8_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_14_b = array_8_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_14_valid_b = array_8_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_15_a = array_8_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_15_valid_a = array_8_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_15_b = array_8_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_15_valid_b = array_8_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_16_a = array_8_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_16_valid_a = array_8_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_16_b = array_8_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_16_valid_b = array_8_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_17_a = array_8_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_17_valid_a = array_8_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_17_b = array_8_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_17_valid_b = array_8_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_18_a = array_8_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_18_valid_a = array_8_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_18_b = array_8_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_18_valid_b = array_8_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_19_a = array_8_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_19_valid_a = array_8_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_19_b = array_8_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_19_valid_b = array_8_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_20_a = array_8_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_20_valid_a = array_8_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_20_b = array_8_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_20_valid_b = array_8_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_21_a = array_8_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_21_valid_a = array_8_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_21_b = array_8_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_21_valid_b = array_8_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_22_a = array_8_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_22_valid_a = array_8_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_22_b = array_8_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_22_valid_b = array_8_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_23_a = array_8_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_23_valid_a = array_8_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_23_b = array_8_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_23_valid_b = array_8_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_24_a = array_8_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_24_valid_a = array_8_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_24_b = array_8_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_24_valid_b = array_8_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_25_a = array_8_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_25_valid_a = array_8_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_25_b = array_8_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_25_valid_b = array_8_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_26_a = array_8_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_26_valid_a = array_8_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_26_b = array_8_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_26_valid_b = array_8_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_27_a = array_8_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_27_valid_a = array_8_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_27_b = array_8_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_27_valid_b = array_8_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_28_a = array_8_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_28_valid_a = array_8_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_28_b = array_8_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_28_valid_b = array_8_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_29_a = array_8_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_29_valid_a = array_8_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_29_b = array_8_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_29_valid_b = array_8_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_30_a = array_8_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_30_valid_a = array_8_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_30_b = array_8_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_30_valid_b = array_8_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_31_a = array_8_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_31_valid_a = array_8_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_9_io_d_in_31_b = array_8_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_9_io_d_in_31_valid_b = array_8_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_9_io_wr_en_mem1 = io_wr_en_mem1_9; // @[BP.scala 325:28]
  assign array_9_io_wr_en_mem2 = io_wr_en_mem2_9; // @[BP.scala 326:28]
  assign array_9_io_wr_en_mem3 = io_wr_en_mem3_9; // @[BP.scala 327:28]
  assign array_9_io_wr_en_mem4 = io_wr_en_mem4_9; // @[BP.scala 328:28]
  assign array_9_io_wr_en_mem5 = io_wr_en_mem5_9; // @[BP.scala 329:28]
  assign array_9_io_wr_en_mem6 = io_wr_en_mem6_9; // @[BP.scala 330:28]
  assign array_9_io_wr_instr_mem1 = io_wr_instr_mem1_9; // @[BP.scala 331:31]
  assign array_9_io_wr_instr_mem2 = io_wr_instr_mem2_9; // @[BP.scala 332:31]
  assign array_9_io_wr_instr_mem3 = io_wr_instr_mem3_9; // @[BP.scala 333:31]
  assign array_9_io_wr_instr_mem4 = io_wr_instr_mem4_9; // @[BP.scala 334:31]
  assign array_9_io_wr_instr_mem5 = io_wr_instr_mem5_9; // @[BP.scala 335:31]
  assign array_9_io_wr_instr_mem6 = io_wr_instr_mem6_9; // @[BP.scala 336:31]
  assign array_9_io_PC1_in = array_8_io_PC6_out; // @[BP.scala 338:24]
  assign array_9_io_Addr_in = array_8_io_Addr_out; // @[BP.scala 339:25]
  assign array_10_clock = clock;
  assign array_10_reset = reset;
  assign array_10_io_d_in_0_a = array_9_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_0_valid_a = array_9_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_0_b = array_9_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_0_valid_b = array_9_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_1_a = array_9_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_1_valid_a = array_9_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_1_b = array_9_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_1_valid_b = array_9_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_2_a = array_9_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_2_valid_a = array_9_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_2_b = array_9_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_2_valid_b = array_9_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_3_a = array_9_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_3_valid_a = array_9_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_3_b = array_9_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_3_valid_b = array_9_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_4_a = array_9_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_4_valid_a = array_9_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_4_b = array_9_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_4_valid_b = array_9_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_5_a = array_9_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_5_valid_a = array_9_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_5_b = array_9_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_5_valid_b = array_9_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_6_a = array_9_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_6_valid_a = array_9_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_6_b = array_9_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_6_valid_b = array_9_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_7_a = array_9_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_7_valid_a = array_9_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_7_b = array_9_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_7_valid_b = array_9_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_8_a = array_9_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_8_valid_a = array_9_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_8_b = array_9_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_8_valid_b = array_9_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_9_a = array_9_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_9_valid_a = array_9_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_9_b = array_9_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_9_valid_b = array_9_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_10_a = array_9_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_10_valid_a = array_9_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_10_b = array_9_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_10_valid_b = array_9_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_11_a = array_9_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_11_valid_a = array_9_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_11_b = array_9_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_11_valid_b = array_9_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_12_a = array_9_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_12_valid_a = array_9_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_12_b = array_9_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_12_valid_b = array_9_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_13_a = array_9_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_13_valid_a = array_9_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_13_b = array_9_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_13_valid_b = array_9_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_14_a = array_9_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_14_valid_a = array_9_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_14_b = array_9_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_14_valid_b = array_9_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_15_a = array_9_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_15_valid_a = array_9_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_15_b = array_9_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_15_valid_b = array_9_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_16_a = array_9_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_16_valid_a = array_9_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_16_b = array_9_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_16_valid_b = array_9_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_17_a = array_9_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_17_valid_a = array_9_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_17_b = array_9_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_17_valid_b = array_9_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_18_a = array_9_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_18_valid_a = array_9_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_18_b = array_9_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_18_valid_b = array_9_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_19_a = array_9_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_19_valid_a = array_9_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_19_b = array_9_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_19_valid_b = array_9_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_20_a = array_9_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_20_valid_a = array_9_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_20_b = array_9_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_20_valid_b = array_9_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_21_a = array_9_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_21_valid_a = array_9_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_21_b = array_9_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_21_valid_b = array_9_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_22_a = array_9_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_22_valid_a = array_9_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_22_b = array_9_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_22_valid_b = array_9_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_23_a = array_9_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_23_valid_a = array_9_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_23_b = array_9_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_23_valid_b = array_9_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_24_a = array_9_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_24_valid_a = array_9_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_24_b = array_9_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_24_valid_b = array_9_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_25_a = array_9_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_25_valid_a = array_9_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_25_b = array_9_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_25_valid_b = array_9_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_26_a = array_9_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_26_valid_a = array_9_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_26_b = array_9_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_26_valid_b = array_9_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_27_a = array_9_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_27_valid_a = array_9_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_27_b = array_9_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_27_valid_b = array_9_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_28_a = array_9_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_28_valid_a = array_9_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_28_b = array_9_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_28_valid_b = array_9_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_29_a = array_9_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_29_valid_a = array_9_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_29_b = array_9_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_29_valid_b = array_9_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_30_a = array_9_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_30_valid_a = array_9_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_30_b = array_9_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_30_valid_b = array_9_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_31_a = array_9_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_31_valid_a = array_9_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_10_io_d_in_31_b = array_9_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_10_io_d_in_31_valid_b = array_9_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_10_io_wr_en_mem1 = io_wr_en_mem1_10; // @[BP.scala 325:28]
  assign array_10_io_wr_en_mem2 = io_wr_en_mem2_10; // @[BP.scala 326:28]
  assign array_10_io_wr_en_mem3 = io_wr_en_mem3_10; // @[BP.scala 327:28]
  assign array_10_io_wr_en_mem4 = io_wr_en_mem4_10; // @[BP.scala 328:28]
  assign array_10_io_wr_en_mem5 = io_wr_en_mem5_10; // @[BP.scala 329:28]
  assign array_10_io_wr_en_mem6 = io_wr_en_mem6_10; // @[BP.scala 330:28]
  assign array_10_io_wr_instr_mem1 = io_wr_instr_mem1_10; // @[BP.scala 331:31]
  assign array_10_io_wr_instr_mem2 = io_wr_instr_mem2_10; // @[BP.scala 332:31]
  assign array_10_io_wr_instr_mem3 = io_wr_instr_mem3_10; // @[BP.scala 333:31]
  assign array_10_io_wr_instr_mem4 = io_wr_instr_mem4_10; // @[BP.scala 334:31]
  assign array_10_io_wr_instr_mem5 = io_wr_instr_mem5_10; // @[BP.scala 335:31]
  assign array_10_io_wr_instr_mem6 = io_wr_instr_mem6_10; // @[BP.scala 336:31]
  assign array_10_io_PC1_in = array_9_io_PC6_out; // @[BP.scala 338:24]
  assign array_10_io_Addr_in = array_9_io_Addr_out; // @[BP.scala 339:25]
  assign array_11_clock = clock;
  assign array_11_reset = reset;
  assign array_11_io_d_in_0_a = array_10_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_0_valid_a = array_10_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_0_b = array_10_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_0_valid_b = array_10_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_1_a = array_10_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_1_valid_a = array_10_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_1_b = array_10_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_1_valid_b = array_10_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_2_a = array_10_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_2_valid_a = array_10_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_2_b = array_10_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_2_valid_b = array_10_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_3_a = array_10_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_3_valid_a = array_10_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_3_b = array_10_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_3_valid_b = array_10_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_4_a = array_10_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_4_valid_a = array_10_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_4_b = array_10_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_4_valid_b = array_10_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_5_a = array_10_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_5_valid_a = array_10_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_5_b = array_10_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_5_valid_b = array_10_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_6_a = array_10_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_6_valid_a = array_10_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_6_b = array_10_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_6_valid_b = array_10_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_7_a = array_10_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_7_valid_a = array_10_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_7_b = array_10_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_7_valid_b = array_10_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_8_a = array_10_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_8_valid_a = array_10_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_8_b = array_10_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_8_valid_b = array_10_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_9_a = array_10_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_9_valid_a = array_10_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_9_b = array_10_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_9_valid_b = array_10_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_10_a = array_10_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_10_valid_a = array_10_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_10_b = array_10_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_10_valid_b = array_10_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_11_a = array_10_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_11_valid_a = array_10_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_11_b = array_10_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_11_valid_b = array_10_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_12_a = array_10_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_12_valid_a = array_10_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_12_b = array_10_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_12_valid_b = array_10_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_13_a = array_10_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_13_valid_a = array_10_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_13_b = array_10_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_13_valid_b = array_10_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_14_a = array_10_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_14_valid_a = array_10_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_14_b = array_10_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_14_valid_b = array_10_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_15_a = array_10_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_15_valid_a = array_10_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_15_b = array_10_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_15_valid_b = array_10_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_16_a = array_10_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_16_valid_a = array_10_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_16_b = array_10_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_16_valid_b = array_10_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_17_a = array_10_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_17_valid_a = array_10_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_17_b = array_10_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_17_valid_b = array_10_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_18_a = array_10_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_18_valid_a = array_10_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_18_b = array_10_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_18_valid_b = array_10_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_19_a = array_10_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_19_valid_a = array_10_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_19_b = array_10_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_19_valid_b = array_10_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_20_a = array_10_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_20_valid_a = array_10_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_20_b = array_10_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_20_valid_b = array_10_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_21_a = array_10_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_21_valid_a = array_10_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_21_b = array_10_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_21_valid_b = array_10_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_22_a = array_10_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_22_valid_a = array_10_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_22_b = array_10_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_22_valid_b = array_10_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_23_a = array_10_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_23_valid_a = array_10_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_23_b = array_10_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_23_valid_b = array_10_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_24_a = array_10_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_24_valid_a = array_10_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_24_b = array_10_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_24_valid_b = array_10_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_25_a = array_10_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_25_valid_a = array_10_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_25_b = array_10_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_25_valid_b = array_10_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_26_a = array_10_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_26_valid_a = array_10_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_26_b = array_10_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_26_valid_b = array_10_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_27_a = array_10_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_27_valid_a = array_10_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_27_b = array_10_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_27_valid_b = array_10_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_28_a = array_10_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_28_valid_a = array_10_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_28_b = array_10_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_28_valid_b = array_10_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_29_a = array_10_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_29_valid_a = array_10_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_29_b = array_10_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_29_valid_b = array_10_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_30_a = array_10_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_30_valid_a = array_10_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_30_b = array_10_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_30_valid_b = array_10_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_31_a = array_10_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_31_valid_a = array_10_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_11_io_d_in_31_b = array_10_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_11_io_d_in_31_valid_b = array_10_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_11_io_wr_en_mem1 = io_wr_en_mem1_11; // @[BP.scala 325:28]
  assign array_11_io_wr_en_mem2 = io_wr_en_mem2_11; // @[BP.scala 326:28]
  assign array_11_io_wr_en_mem3 = io_wr_en_mem3_11; // @[BP.scala 327:28]
  assign array_11_io_wr_en_mem4 = io_wr_en_mem4_11; // @[BP.scala 328:28]
  assign array_11_io_wr_en_mem5 = io_wr_en_mem5_11; // @[BP.scala 329:28]
  assign array_11_io_wr_en_mem6 = io_wr_en_mem6_11; // @[BP.scala 330:28]
  assign array_11_io_wr_instr_mem1 = io_wr_instr_mem1_11; // @[BP.scala 331:31]
  assign array_11_io_wr_instr_mem2 = io_wr_instr_mem2_11; // @[BP.scala 332:31]
  assign array_11_io_wr_instr_mem3 = io_wr_instr_mem3_11; // @[BP.scala 333:31]
  assign array_11_io_wr_instr_mem4 = io_wr_instr_mem4_11; // @[BP.scala 334:31]
  assign array_11_io_wr_instr_mem5 = io_wr_instr_mem5_11; // @[BP.scala 335:31]
  assign array_11_io_wr_instr_mem6 = io_wr_instr_mem6_11; // @[BP.scala 336:31]
  assign array_11_io_PC1_in = array_10_io_PC6_out; // @[BP.scala 338:24]
  assign array_11_io_Addr_in = array_10_io_Addr_out; // @[BP.scala 339:25]
  assign array_12_clock = clock;
  assign array_12_reset = reset;
  assign array_12_io_d_in_0_a = array_11_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_0_valid_a = array_11_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_0_b = array_11_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_0_valid_b = array_11_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_1_a = array_11_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_1_valid_a = array_11_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_1_b = array_11_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_1_valid_b = array_11_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_2_a = array_11_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_2_valid_a = array_11_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_2_b = array_11_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_2_valid_b = array_11_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_3_a = array_11_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_3_valid_a = array_11_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_3_b = array_11_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_3_valid_b = array_11_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_4_a = array_11_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_4_valid_a = array_11_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_4_b = array_11_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_4_valid_b = array_11_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_5_a = array_11_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_5_valid_a = array_11_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_5_b = array_11_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_5_valid_b = array_11_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_6_a = array_11_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_6_valid_a = array_11_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_6_b = array_11_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_6_valid_b = array_11_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_7_a = array_11_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_7_valid_a = array_11_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_7_b = array_11_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_7_valid_b = array_11_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_8_a = array_11_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_8_valid_a = array_11_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_8_b = array_11_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_8_valid_b = array_11_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_9_a = array_11_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_9_valid_a = array_11_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_9_b = array_11_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_9_valid_b = array_11_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_10_a = array_11_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_10_valid_a = array_11_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_10_b = array_11_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_10_valid_b = array_11_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_11_a = array_11_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_11_valid_a = array_11_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_11_b = array_11_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_11_valid_b = array_11_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_12_a = array_11_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_12_valid_a = array_11_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_12_b = array_11_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_12_valid_b = array_11_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_13_a = array_11_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_13_valid_a = array_11_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_13_b = array_11_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_13_valid_b = array_11_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_14_a = array_11_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_14_valid_a = array_11_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_14_b = array_11_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_14_valid_b = array_11_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_15_a = array_11_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_15_valid_a = array_11_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_15_b = array_11_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_15_valid_b = array_11_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_16_a = array_11_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_16_valid_a = array_11_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_16_b = array_11_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_16_valid_b = array_11_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_17_a = array_11_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_17_valid_a = array_11_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_17_b = array_11_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_17_valid_b = array_11_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_18_a = array_11_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_18_valid_a = array_11_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_18_b = array_11_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_18_valid_b = array_11_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_19_a = array_11_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_19_valid_a = array_11_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_19_b = array_11_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_19_valid_b = array_11_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_20_a = array_11_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_20_valid_a = array_11_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_20_b = array_11_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_20_valid_b = array_11_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_21_a = array_11_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_21_valid_a = array_11_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_21_b = array_11_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_21_valid_b = array_11_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_22_a = array_11_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_22_valid_a = array_11_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_22_b = array_11_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_22_valid_b = array_11_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_23_a = array_11_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_23_valid_a = array_11_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_23_b = array_11_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_23_valid_b = array_11_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_24_a = array_11_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_24_valid_a = array_11_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_24_b = array_11_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_24_valid_b = array_11_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_25_a = array_11_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_25_valid_a = array_11_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_25_b = array_11_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_25_valid_b = array_11_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_26_a = array_11_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_26_valid_a = array_11_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_26_b = array_11_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_26_valid_b = array_11_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_27_a = array_11_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_27_valid_a = array_11_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_27_b = array_11_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_27_valid_b = array_11_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_28_a = array_11_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_28_valid_a = array_11_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_28_b = array_11_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_28_valid_b = array_11_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_29_a = array_11_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_29_valid_a = array_11_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_29_b = array_11_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_29_valid_b = array_11_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_30_a = array_11_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_30_valid_a = array_11_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_30_b = array_11_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_30_valid_b = array_11_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_31_a = array_11_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_31_valid_a = array_11_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_12_io_d_in_31_b = array_11_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_12_io_d_in_31_valid_b = array_11_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_12_io_wr_en_mem1 = io_wr_en_mem1_12; // @[BP.scala 325:28]
  assign array_12_io_wr_en_mem2 = io_wr_en_mem2_12; // @[BP.scala 326:28]
  assign array_12_io_wr_en_mem3 = io_wr_en_mem3_12; // @[BP.scala 327:28]
  assign array_12_io_wr_en_mem4 = io_wr_en_mem4_12; // @[BP.scala 328:28]
  assign array_12_io_wr_en_mem5 = io_wr_en_mem5_12; // @[BP.scala 329:28]
  assign array_12_io_wr_en_mem6 = io_wr_en_mem6_12; // @[BP.scala 330:28]
  assign array_12_io_wr_instr_mem1 = io_wr_instr_mem1_12; // @[BP.scala 331:31]
  assign array_12_io_wr_instr_mem2 = io_wr_instr_mem2_12; // @[BP.scala 332:31]
  assign array_12_io_wr_instr_mem3 = io_wr_instr_mem3_12; // @[BP.scala 333:31]
  assign array_12_io_wr_instr_mem4 = io_wr_instr_mem4_12; // @[BP.scala 334:31]
  assign array_12_io_wr_instr_mem5 = io_wr_instr_mem5_12; // @[BP.scala 335:31]
  assign array_12_io_wr_instr_mem6 = io_wr_instr_mem6_12; // @[BP.scala 336:31]
  assign array_12_io_PC1_in = array_11_io_PC6_out; // @[BP.scala 338:24]
  assign array_12_io_Addr_in = array_11_io_Addr_out; // @[BP.scala 339:25]
  assign array_13_clock = clock;
  assign array_13_reset = reset;
  assign array_13_io_d_in_0_a = array_12_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_0_valid_a = array_12_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_0_b = array_12_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_0_valid_b = array_12_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_1_a = array_12_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_1_valid_a = array_12_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_1_b = array_12_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_1_valid_b = array_12_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_2_a = array_12_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_2_valid_a = array_12_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_2_b = array_12_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_2_valid_b = array_12_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_3_a = array_12_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_3_valid_a = array_12_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_3_b = array_12_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_3_valid_b = array_12_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_4_a = array_12_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_4_valid_a = array_12_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_4_b = array_12_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_4_valid_b = array_12_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_5_a = array_12_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_5_valid_a = array_12_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_5_b = array_12_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_5_valid_b = array_12_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_6_a = array_12_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_6_valid_a = array_12_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_6_b = array_12_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_6_valid_b = array_12_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_7_a = array_12_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_7_valid_a = array_12_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_7_b = array_12_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_7_valid_b = array_12_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_8_a = array_12_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_8_valid_a = array_12_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_8_b = array_12_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_8_valid_b = array_12_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_9_a = array_12_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_9_valid_a = array_12_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_9_b = array_12_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_9_valid_b = array_12_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_10_a = array_12_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_10_valid_a = array_12_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_10_b = array_12_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_10_valid_b = array_12_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_11_a = array_12_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_11_valid_a = array_12_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_11_b = array_12_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_11_valid_b = array_12_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_12_a = array_12_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_12_valid_a = array_12_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_12_b = array_12_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_12_valid_b = array_12_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_13_a = array_12_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_13_valid_a = array_12_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_13_b = array_12_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_13_valid_b = array_12_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_14_a = array_12_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_14_valid_a = array_12_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_14_b = array_12_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_14_valid_b = array_12_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_15_a = array_12_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_15_valid_a = array_12_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_15_b = array_12_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_15_valid_b = array_12_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_16_a = array_12_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_16_valid_a = array_12_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_16_b = array_12_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_16_valid_b = array_12_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_17_a = array_12_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_17_valid_a = array_12_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_17_b = array_12_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_17_valid_b = array_12_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_18_a = array_12_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_18_valid_a = array_12_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_18_b = array_12_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_18_valid_b = array_12_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_19_a = array_12_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_19_valid_a = array_12_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_19_b = array_12_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_19_valid_b = array_12_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_20_a = array_12_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_20_valid_a = array_12_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_20_b = array_12_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_20_valid_b = array_12_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_21_a = array_12_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_21_valid_a = array_12_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_21_b = array_12_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_21_valid_b = array_12_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_22_a = array_12_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_22_valid_a = array_12_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_22_b = array_12_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_22_valid_b = array_12_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_23_a = array_12_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_23_valid_a = array_12_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_23_b = array_12_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_23_valid_b = array_12_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_24_a = array_12_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_24_valid_a = array_12_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_24_b = array_12_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_24_valid_b = array_12_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_25_a = array_12_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_25_valid_a = array_12_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_25_b = array_12_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_25_valid_b = array_12_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_26_a = array_12_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_26_valid_a = array_12_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_26_b = array_12_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_26_valid_b = array_12_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_27_a = array_12_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_27_valid_a = array_12_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_27_b = array_12_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_27_valid_b = array_12_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_28_a = array_12_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_28_valid_a = array_12_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_28_b = array_12_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_28_valid_b = array_12_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_29_a = array_12_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_29_valid_a = array_12_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_29_b = array_12_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_29_valid_b = array_12_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_30_a = array_12_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_30_valid_a = array_12_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_30_b = array_12_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_30_valid_b = array_12_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_31_a = array_12_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_31_valid_a = array_12_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_13_io_d_in_31_b = array_12_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_13_io_d_in_31_valid_b = array_12_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_13_io_wr_en_mem1 = io_wr_en_mem1_13; // @[BP.scala 325:28]
  assign array_13_io_wr_en_mem2 = io_wr_en_mem2_13; // @[BP.scala 326:28]
  assign array_13_io_wr_en_mem3 = io_wr_en_mem3_13; // @[BP.scala 327:28]
  assign array_13_io_wr_en_mem4 = io_wr_en_mem4_13; // @[BP.scala 328:28]
  assign array_13_io_wr_en_mem5 = io_wr_en_mem5_13; // @[BP.scala 329:28]
  assign array_13_io_wr_en_mem6 = io_wr_en_mem6_13; // @[BP.scala 330:28]
  assign array_13_io_wr_instr_mem1 = io_wr_instr_mem1_13; // @[BP.scala 331:31]
  assign array_13_io_wr_instr_mem2 = io_wr_instr_mem2_13; // @[BP.scala 332:31]
  assign array_13_io_wr_instr_mem3 = io_wr_instr_mem3_13; // @[BP.scala 333:31]
  assign array_13_io_wr_instr_mem4 = io_wr_instr_mem4_13; // @[BP.scala 334:31]
  assign array_13_io_wr_instr_mem5 = io_wr_instr_mem5_13; // @[BP.scala 335:31]
  assign array_13_io_wr_instr_mem6 = io_wr_instr_mem6_13; // @[BP.scala 336:31]
  assign array_13_io_PC1_in = array_12_io_PC6_out; // @[BP.scala 338:24]
  assign array_13_io_Addr_in = array_12_io_Addr_out; // @[BP.scala 339:25]
  assign array_14_clock = clock;
  assign array_14_reset = reset;
  assign array_14_io_d_in_0_a = array_13_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_0_valid_a = array_13_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_0_b = array_13_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_0_valid_b = array_13_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_1_a = array_13_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_1_valid_a = array_13_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_1_b = array_13_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_1_valid_b = array_13_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_2_a = array_13_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_2_valid_a = array_13_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_2_b = array_13_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_2_valid_b = array_13_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_3_a = array_13_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_3_valid_a = array_13_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_3_b = array_13_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_3_valid_b = array_13_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_4_a = array_13_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_4_valid_a = array_13_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_4_b = array_13_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_4_valid_b = array_13_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_5_a = array_13_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_5_valid_a = array_13_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_5_b = array_13_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_5_valid_b = array_13_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_6_a = array_13_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_6_valid_a = array_13_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_6_b = array_13_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_6_valid_b = array_13_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_7_a = array_13_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_7_valid_a = array_13_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_7_b = array_13_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_7_valid_b = array_13_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_8_a = array_13_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_8_valid_a = array_13_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_8_b = array_13_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_8_valid_b = array_13_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_9_a = array_13_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_9_valid_a = array_13_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_9_b = array_13_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_9_valid_b = array_13_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_10_a = array_13_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_10_valid_a = array_13_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_10_b = array_13_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_10_valid_b = array_13_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_11_a = array_13_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_11_valid_a = array_13_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_11_b = array_13_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_11_valid_b = array_13_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_12_a = array_13_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_12_valid_a = array_13_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_12_b = array_13_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_12_valid_b = array_13_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_13_a = array_13_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_13_valid_a = array_13_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_13_b = array_13_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_13_valid_b = array_13_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_14_a = array_13_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_14_valid_a = array_13_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_14_b = array_13_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_14_valid_b = array_13_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_15_a = array_13_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_15_valid_a = array_13_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_15_b = array_13_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_15_valid_b = array_13_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_16_a = array_13_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_16_valid_a = array_13_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_16_b = array_13_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_16_valid_b = array_13_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_17_a = array_13_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_17_valid_a = array_13_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_17_b = array_13_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_17_valid_b = array_13_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_18_a = array_13_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_18_valid_a = array_13_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_18_b = array_13_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_18_valid_b = array_13_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_19_a = array_13_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_19_valid_a = array_13_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_19_b = array_13_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_19_valid_b = array_13_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_20_a = array_13_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_20_valid_a = array_13_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_20_b = array_13_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_20_valid_b = array_13_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_21_a = array_13_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_21_valid_a = array_13_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_21_b = array_13_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_21_valid_b = array_13_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_22_a = array_13_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_22_valid_a = array_13_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_22_b = array_13_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_22_valid_b = array_13_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_23_a = array_13_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_23_valid_a = array_13_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_23_b = array_13_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_23_valid_b = array_13_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_24_a = array_13_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_24_valid_a = array_13_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_24_b = array_13_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_24_valid_b = array_13_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_25_a = array_13_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_25_valid_a = array_13_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_25_b = array_13_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_25_valid_b = array_13_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_26_a = array_13_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_26_valid_a = array_13_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_26_b = array_13_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_26_valid_b = array_13_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_27_a = array_13_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_27_valid_a = array_13_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_27_b = array_13_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_27_valid_b = array_13_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_28_a = array_13_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_28_valid_a = array_13_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_28_b = array_13_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_28_valid_b = array_13_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_29_a = array_13_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_29_valid_a = array_13_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_29_b = array_13_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_29_valid_b = array_13_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_30_a = array_13_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_30_valid_a = array_13_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_30_b = array_13_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_30_valid_b = array_13_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_31_a = array_13_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_31_valid_a = array_13_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_14_io_d_in_31_b = array_13_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_14_io_d_in_31_valid_b = array_13_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_14_io_wr_en_mem1 = io_wr_en_mem1_14; // @[BP.scala 325:28]
  assign array_14_io_wr_en_mem2 = io_wr_en_mem2_14; // @[BP.scala 326:28]
  assign array_14_io_wr_en_mem3 = io_wr_en_mem3_14; // @[BP.scala 327:28]
  assign array_14_io_wr_en_mem4 = io_wr_en_mem4_14; // @[BP.scala 328:28]
  assign array_14_io_wr_en_mem5 = io_wr_en_mem5_14; // @[BP.scala 329:28]
  assign array_14_io_wr_en_mem6 = io_wr_en_mem6_14; // @[BP.scala 330:28]
  assign array_14_io_wr_instr_mem1 = io_wr_instr_mem1_14; // @[BP.scala 331:31]
  assign array_14_io_wr_instr_mem2 = io_wr_instr_mem2_14; // @[BP.scala 332:31]
  assign array_14_io_wr_instr_mem3 = io_wr_instr_mem3_14; // @[BP.scala 333:31]
  assign array_14_io_wr_instr_mem4 = io_wr_instr_mem4_14; // @[BP.scala 334:31]
  assign array_14_io_wr_instr_mem5 = io_wr_instr_mem5_14; // @[BP.scala 335:31]
  assign array_14_io_wr_instr_mem6 = io_wr_instr_mem6_14; // @[BP.scala 336:31]
  assign array_14_io_PC1_in = array_13_io_PC6_out; // @[BP.scala 338:24]
  assign array_14_io_Addr_in = array_13_io_Addr_out; // @[BP.scala 339:25]
  assign array_15_clock = clock;
  assign array_15_reset = reset;
  assign array_15_io_d_in_0_a = array_14_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_0_valid_a = array_14_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_0_b = array_14_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_0_valid_b = array_14_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_1_a = array_14_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_1_valid_a = array_14_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_1_b = array_14_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_1_valid_b = array_14_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_2_a = array_14_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_2_valid_a = array_14_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_2_b = array_14_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_2_valid_b = array_14_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_3_a = array_14_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_3_valid_a = array_14_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_3_b = array_14_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_3_valid_b = array_14_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_4_a = array_14_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_4_valid_a = array_14_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_4_b = array_14_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_4_valid_b = array_14_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_5_a = array_14_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_5_valid_a = array_14_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_5_b = array_14_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_5_valid_b = array_14_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_6_a = array_14_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_6_valid_a = array_14_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_6_b = array_14_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_6_valid_b = array_14_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_7_a = array_14_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_7_valid_a = array_14_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_7_b = array_14_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_7_valid_b = array_14_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_8_a = array_14_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_8_valid_a = array_14_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_8_b = array_14_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_8_valid_b = array_14_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_9_a = array_14_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_9_valid_a = array_14_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_9_b = array_14_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_9_valid_b = array_14_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_10_a = array_14_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_10_valid_a = array_14_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_10_b = array_14_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_10_valid_b = array_14_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_11_a = array_14_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_11_valid_a = array_14_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_11_b = array_14_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_11_valid_b = array_14_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_12_a = array_14_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_12_valid_a = array_14_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_12_b = array_14_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_12_valid_b = array_14_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_13_a = array_14_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_13_valid_a = array_14_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_13_b = array_14_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_13_valid_b = array_14_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_14_a = array_14_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_14_valid_a = array_14_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_14_b = array_14_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_14_valid_b = array_14_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_15_a = array_14_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_15_valid_a = array_14_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_15_b = array_14_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_15_valid_b = array_14_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_16_a = array_14_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_16_valid_a = array_14_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_16_b = array_14_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_16_valid_b = array_14_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_17_a = array_14_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_17_valid_a = array_14_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_17_b = array_14_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_17_valid_b = array_14_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_18_a = array_14_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_18_valid_a = array_14_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_18_b = array_14_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_18_valid_b = array_14_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_19_a = array_14_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_19_valid_a = array_14_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_19_b = array_14_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_19_valid_b = array_14_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_20_a = array_14_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_20_valid_a = array_14_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_20_b = array_14_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_20_valid_b = array_14_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_21_a = array_14_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_21_valid_a = array_14_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_21_b = array_14_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_21_valid_b = array_14_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_22_a = array_14_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_22_valid_a = array_14_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_22_b = array_14_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_22_valid_b = array_14_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_23_a = array_14_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_23_valid_a = array_14_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_23_b = array_14_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_23_valid_b = array_14_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_24_a = array_14_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_24_valid_a = array_14_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_24_b = array_14_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_24_valid_b = array_14_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_25_a = array_14_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_25_valid_a = array_14_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_25_b = array_14_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_25_valid_b = array_14_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_26_a = array_14_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_26_valid_a = array_14_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_26_b = array_14_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_26_valid_b = array_14_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_27_a = array_14_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_27_valid_a = array_14_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_27_b = array_14_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_27_valid_b = array_14_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_28_a = array_14_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_28_valid_a = array_14_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_28_b = array_14_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_28_valid_b = array_14_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_29_a = array_14_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_29_valid_a = array_14_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_29_b = array_14_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_29_valid_b = array_14_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_30_a = array_14_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_30_valid_a = array_14_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_30_b = array_14_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_30_valid_b = array_14_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_31_a = array_14_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_31_valid_a = array_14_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_15_io_d_in_31_b = array_14_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_15_io_d_in_31_valid_b = array_14_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_15_io_wr_en_mem1 = io_wr_en_mem1_15; // @[BP.scala 325:28]
  assign array_15_io_wr_en_mem2 = io_wr_en_mem2_15; // @[BP.scala 326:28]
  assign array_15_io_wr_en_mem3 = io_wr_en_mem3_15; // @[BP.scala 327:28]
  assign array_15_io_wr_en_mem4 = io_wr_en_mem4_15; // @[BP.scala 328:28]
  assign array_15_io_wr_en_mem5 = io_wr_en_mem5_15; // @[BP.scala 329:28]
  assign array_15_io_wr_en_mem6 = io_wr_en_mem6_15; // @[BP.scala 330:28]
  assign array_15_io_wr_instr_mem1 = io_wr_instr_mem1_15; // @[BP.scala 331:31]
  assign array_15_io_wr_instr_mem2 = io_wr_instr_mem2_15; // @[BP.scala 332:31]
  assign array_15_io_wr_instr_mem3 = io_wr_instr_mem3_15; // @[BP.scala 333:31]
  assign array_15_io_wr_instr_mem4 = io_wr_instr_mem4_15; // @[BP.scala 334:31]
  assign array_15_io_wr_instr_mem5 = io_wr_instr_mem5_15; // @[BP.scala 335:31]
  assign array_15_io_wr_instr_mem6 = io_wr_instr_mem6_15; // @[BP.scala 336:31]
  assign array_15_io_PC1_in = array_14_io_PC6_out; // @[BP.scala 338:24]
  assign array_15_io_Addr_in = array_14_io_Addr_out; // @[BP.scala 339:25]
  assign array_16_clock = clock;
  assign array_16_reset = reset;
  assign array_16_io_d_in_0_a = array_15_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_0_valid_a = array_15_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_0_b = array_15_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_0_valid_b = array_15_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_1_a = array_15_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_1_valid_a = array_15_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_1_b = array_15_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_1_valid_b = array_15_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_2_a = array_15_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_2_valid_a = array_15_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_2_b = array_15_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_2_valid_b = array_15_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_3_a = array_15_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_3_valid_a = array_15_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_3_b = array_15_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_3_valid_b = array_15_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_4_a = array_15_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_4_valid_a = array_15_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_4_b = array_15_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_4_valid_b = array_15_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_5_a = array_15_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_5_valid_a = array_15_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_5_b = array_15_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_5_valid_b = array_15_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_6_a = array_15_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_6_valid_a = array_15_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_6_b = array_15_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_6_valid_b = array_15_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_7_a = array_15_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_7_valid_a = array_15_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_7_b = array_15_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_7_valid_b = array_15_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_8_a = array_15_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_8_valid_a = array_15_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_8_b = array_15_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_8_valid_b = array_15_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_9_a = array_15_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_9_valid_a = array_15_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_9_b = array_15_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_9_valid_b = array_15_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_10_a = array_15_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_10_valid_a = array_15_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_10_b = array_15_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_10_valid_b = array_15_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_11_a = array_15_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_11_valid_a = array_15_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_11_b = array_15_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_11_valid_b = array_15_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_12_a = array_15_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_12_valid_a = array_15_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_12_b = array_15_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_12_valid_b = array_15_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_13_a = array_15_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_13_valid_a = array_15_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_13_b = array_15_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_13_valid_b = array_15_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_14_a = array_15_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_14_valid_a = array_15_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_14_b = array_15_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_14_valid_b = array_15_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_15_a = array_15_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_15_valid_a = array_15_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_15_b = array_15_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_15_valid_b = array_15_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_16_a = array_15_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_16_valid_a = array_15_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_16_b = array_15_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_16_valid_b = array_15_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_17_a = array_15_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_17_valid_a = array_15_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_17_b = array_15_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_17_valid_b = array_15_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_18_a = array_15_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_18_valid_a = array_15_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_18_b = array_15_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_18_valid_b = array_15_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_19_a = array_15_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_19_valid_a = array_15_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_19_b = array_15_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_19_valid_b = array_15_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_20_a = array_15_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_20_valid_a = array_15_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_20_b = array_15_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_20_valid_b = array_15_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_21_a = array_15_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_21_valid_a = array_15_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_21_b = array_15_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_21_valid_b = array_15_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_22_a = array_15_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_22_valid_a = array_15_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_22_b = array_15_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_22_valid_b = array_15_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_23_a = array_15_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_23_valid_a = array_15_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_23_b = array_15_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_23_valid_b = array_15_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_24_a = array_15_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_24_valid_a = array_15_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_24_b = array_15_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_24_valid_b = array_15_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_25_a = array_15_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_25_valid_a = array_15_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_25_b = array_15_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_25_valid_b = array_15_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_26_a = array_15_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_26_valid_a = array_15_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_26_b = array_15_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_26_valid_b = array_15_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_27_a = array_15_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_27_valid_a = array_15_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_27_b = array_15_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_27_valid_b = array_15_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_28_a = array_15_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_28_valid_a = array_15_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_28_b = array_15_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_28_valid_b = array_15_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_29_a = array_15_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_29_valid_a = array_15_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_29_b = array_15_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_29_valid_b = array_15_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_30_a = array_15_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_30_valid_a = array_15_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_30_b = array_15_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_30_valid_b = array_15_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_31_a = array_15_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_31_valid_a = array_15_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_16_io_d_in_31_b = array_15_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_16_io_d_in_31_valid_b = array_15_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_16_io_wr_en_mem1 = io_wr_en_mem1_16; // @[BP.scala 325:28]
  assign array_16_io_wr_en_mem2 = io_wr_en_mem2_16; // @[BP.scala 326:28]
  assign array_16_io_wr_en_mem3 = io_wr_en_mem3_16; // @[BP.scala 327:28]
  assign array_16_io_wr_en_mem4 = io_wr_en_mem4_16; // @[BP.scala 328:28]
  assign array_16_io_wr_en_mem5 = io_wr_en_mem5_16; // @[BP.scala 329:28]
  assign array_16_io_wr_en_mem6 = io_wr_en_mem6_16; // @[BP.scala 330:28]
  assign array_16_io_wr_instr_mem1 = io_wr_instr_mem1_16; // @[BP.scala 331:31]
  assign array_16_io_wr_instr_mem2 = io_wr_instr_mem2_16; // @[BP.scala 332:31]
  assign array_16_io_wr_instr_mem3 = io_wr_instr_mem3_16; // @[BP.scala 333:31]
  assign array_16_io_wr_instr_mem4 = io_wr_instr_mem4_16; // @[BP.scala 334:31]
  assign array_16_io_wr_instr_mem5 = io_wr_instr_mem5_16; // @[BP.scala 335:31]
  assign array_16_io_wr_instr_mem6 = io_wr_instr_mem6_16; // @[BP.scala 336:31]
  assign array_16_io_PC1_in = array_15_io_PC6_out; // @[BP.scala 338:24]
  assign array_16_io_Addr_in = array_15_io_Addr_out; // @[BP.scala 339:25]
  assign array_17_clock = clock;
  assign array_17_reset = reset;
  assign array_17_io_d_in_0_a = array_16_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_0_valid_a = array_16_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_0_b = array_16_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_0_valid_b = array_16_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_1_a = array_16_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_1_valid_a = array_16_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_1_b = array_16_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_1_valid_b = array_16_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_2_a = array_16_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_2_valid_a = array_16_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_2_b = array_16_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_2_valid_b = array_16_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_3_a = array_16_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_3_valid_a = array_16_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_3_b = array_16_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_3_valid_b = array_16_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_4_a = array_16_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_4_valid_a = array_16_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_4_b = array_16_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_4_valid_b = array_16_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_5_a = array_16_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_5_valid_a = array_16_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_5_b = array_16_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_5_valid_b = array_16_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_6_a = array_16_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_6_valid_a = array_16_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_6_b = array_16_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_6_valid_b = array_16_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_7_a = array_16_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_7_valid_a = array_16_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_7_b = array_16_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_7_valid_b = array_16_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_8_a = array_16_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_8_valid_a = array_16_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_8_b = array_16_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_8_valid_b = array_16_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_9_a = array_16_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_9_valid_a = array_16_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_9_b = array_16_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_9_valid_b = array_16_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_10_a = array_16_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_10_valid_a = array_16_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_10_b = array_16_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_10_valid_b = array_16_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_11_a = array_16_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_11_valid_a = array_16_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_11_b = array_16_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_11_valid_b = array_16_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_12_a = array_16_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_12_valid_a = array_16_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_12_b = array_16_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_12_valid_b = array_16_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_13_a = array_16_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_13_valid_a = array_16_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_13_b = array_16_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_13_valid_b = array_16_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_14_a = array_16_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_14_valid_a = array_16_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_14_b = array_16_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_14_valid_b = array_16_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_15_a = array_16_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_15_valid_a = array_16_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_15_b = array_16_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_15_valid_b = array_16_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_16_a = array_16_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_16_valid_a = array_16_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_16_b = array_16_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_16_valid_b = array_16_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_17_a = array_16_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_17_valid_a = array_16_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_17_b = array_16_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_17_valid_b = array_16_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_18_a = array_16_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_18_valid_a = array_16_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_18_b = array_16_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_18_valid_b = array_16_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_19_a = array_16_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_19_valid_a = array_16_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_19_b = array_16_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_19_valid_b = array_16_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_20_a = array_16_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_20_valid_a = array_16_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_20_b = array_16_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_20_valid_b = array_16_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_21_a = array_16_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_21_valid_a = array_16_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_21_b = array_16_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_21_valid_b = array_16_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_22_a = array_16_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_22_valid_a = array_16_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_22_b = array_16_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_22_valid_b = array_16_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_23_a = array_16_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_23_valid_a = array_16_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_23_b = array_16_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_23_valid_b = array_16_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_24_a = array_16_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_24_valid_a = array_16_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_24_b = array_16_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_24_valid_b = array_16_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_25_a = array_16_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_25_valid_a = array_16_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_25_b = array_16_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_25_valid_b = array_16_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_26_a = array_16_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_26_valid_a = array_16_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_26_b = array_16_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_26_valid_b = array_16_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_27_a = array_16_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_27_valid_a = array_16_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_27_b = array_16_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_27_valid_b = array_16_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_28_a = array_16_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_28_valid_a = array_16_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_28_b = array_16_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_28_valid_b = array_16_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_29_a = array_16_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_29_valid_a = array_16_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_29_b = array_16_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_29_valid_b = array_16_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_30_a = array_16_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_30_valid_a = array_16_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_30_b = array_16_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_30_valid_b = array_16_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_31_a = array_16_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_31_valid_a = array_16_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_17_io_d_in_31_b = array_16_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_17_io_d_in_31_valid_b = array_16_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_17_io_wr_en_mem1 = io_wr_en_mem1_17; // @[BP.scala 325:28]
  assign array_17_io_wr_en_mem2 = io_wr_en_mem2_17; // @[BP.scala 326:28]
  assign array_17_io_wr_en_mem3 = io_wr_en_mem3_17; // @[BP.scala 327:28]
  assign array_17_io_wr_en_mem4 = io_wr_en_mem4_17; // @[BP.scala 328:28]
  assign array_17_io_wr_en_mem5 = io_wr_en_mem5_17; // @[BP.scala 329:28]
  assign array_17_io_wr_en_mem6 = io_wr_en_mem6_17; // @[BP.scala 330:28]
  assign array_17_io_wr_instr_mem1 = io_wr_instr_mem1_17; // @[BP.scala 331:31]
  assign array_17_io_wr_instr_mem2 = io_wr_instr_mem2_17; // @[BP.scala 332:31]
  assign array_17_io_wr_instr_mem3 = io_wr_instr_mem3_17; // @[BP.scala 333:31]
  assign array_17_io_wr_instr_mem4 = io_wr_instr_mem4_17; // @[BP.scala 334:31]
  assign array_17_io_wr_instr_mem5 = io_wr_instr_mem5_17; // @[BP.scala 335:31]
  assign array_17_io_wr_instr_mem6 = io_wr_instr_mem6_17; // @[BP.scala 336:31]
  assign array_17_io_PC1_in = array_16_io_PC6_out; // @[BP.scala 338:24]
  assign array_17_io_Addr_in = array_16_io_Addr_out; // @[BP.scala 339:25]
  assign array_18_clock = clock;
  assign array_18_reset = reset;
  assign array_18_io_d_in_0_a = array_17_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_0_valid_a = array_17_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_0_b = array_17_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_0_valid_b = array_17_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_1_a = array_17_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_1_valid_a = array_17_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_1_b = array_17_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_1_valid_b = array_17_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_2_a = array_17_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_2_valid_a = array_17_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_2_b = array_17_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_2_valid_b = array_17_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_3_a = array_17_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_3_valid_a = array_17_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_3_b = array_17_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_3_valid_b = array_17_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_4_a = array_17_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_4_valid_a = array_17_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_4_b = array_17_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_4_valid_b = array_17_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_5_a = array_17_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_5_valid_a = array_17_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_5_b = array_17_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_5_valid_b = array_17_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_6_a = array_17_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_6_valid_a = array_17_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_6_b = array_17_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_6_valid_b = array_17_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_7_a = array_17_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_7_valid_a = array_17_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_7_b = array_17_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_7_valid_b = array_17_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_8_a = array_17_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_8_valid_a = array_17_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_8_b = array_17_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_8_valid_b = array_17_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_9_a = array_17_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_9_valid_a = array_17_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_9_b = array_17_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_9_valid_b = array_17_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_10_a = array_17_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_10_valid_a = array_17_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_10_b = array_17_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_10_valid_b = array_17_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_11_a = array_17_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_11_valid_a = array_17_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_11_b = array_17_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_11_valid_b = array_17_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_12_a = array_17_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_12_valid_a = array_17_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_12_b = array_17_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_12_valid_b = array_17_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_13_a = array_17_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_13_valid_a = array_17_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_13_b = array_17_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_13_valid_b = array_17_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_14_a = array_17_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_14_valid_a = array_17_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_14_b = array_17_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_14_valid_b = array_17_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_15_a = array_17_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_15_valid_a = array_17_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_15_b = array_17_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_15_valid_b = array_17_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_16_a = array_17_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_16_valid_a = array_17_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_16_b = array_17_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_16_valid_b = array_17_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_17_a = array_17_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_17_valid_a = array_17_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_17_b = array_17_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_17_valid_b = array_17_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_18_a = array_17_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_18_valid_a = array_17_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_18_b = array_17_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_18_valid_b = array_17_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_19_a = array_17_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_19_valid_a = array_17_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_19_b = array_17_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_19_valid_b = array_17_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_20_a = array_17_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_20_valid_a = array_17_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_20_b = array_17_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_20_valid_b = array_17_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_21_a = array_17_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_21_valid_a = array_17_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_21_b = array_17_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_21_valid_b = array_17_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_22_a = array_17_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_22_valid_a = array_17_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_22_b = array_17_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_22_valid_b = array_17_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_23_a = array_17_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_23_valid_a = array_17_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_23_b = array_17_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_23_valid_b = array_17_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_24_a = array_17_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_24_valid_a = array_17_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_24_b = array_17_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_24_valid_b = array_17_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_25_a = array_17_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_25_valid_a = array_17_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_25_b = array_17_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_25_valid_b = array_17_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_26_a = array_17_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_26_valid_a = array_17_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_26_b = array_17_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_26_valid_b = array_17_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_27_a = array_17_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_27_valid_a = array_17_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_27_b = array_17_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_27_valid_b = array_17_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_28_a = array_17_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_28_valid_a = array_17_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_28_b = array_17_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_28_valid_b = array_17_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_29_a = array_17_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_29_valid_a = array_17_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_29_b = array_17_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_29_valid_b = array_17_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_30_a = array_17_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_30_valid_a = array_17_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_30_b = array_17_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_30_valid_b = array_17_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_31_a = array_17_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_31_valid_a = array_17_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_18_io_d_in_31_b = array_17_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_18_io_d_in_31_valid_b = array_17_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_18_io_wr_en_mem1 = io_wr_en_mem1_18; // @[BP.scala 325:28]
  assign array_18_io_wr_en_mem2 = io_wr_en_mem2_18; // @[BP.scala 326:28]
  assign array_18_io_wr_en_mem3 = io_wr_en_mem3_18; // @[BP.scala 327:28]
  assign array_18_io_wr_en_mem4 = io_wr_en_mem4_18; // @[BP.scala 328:28]
  assign array_18_io_wr_en_mem5 = io_wr_en_mem5_18; // @[BP.scala 329:28]
  assign array_18_io_wr_en_mem6 = io_wr_en_mem6_18; // @[BP.scala 330:28]
  assign array_18_io_wr_instr_mem1 = io_wr_instr_mem1_18; // @[BP.scala 331:31]
  assign array_18_io_wr_instr_mem2 = io_wr_instr_mem2_18; // @[BP.scala 332:31]
  assign array_18_io_wr_instr_mem3 = io_wr_instr_mem3_18; // @[BP.scala 333:31]
  assign array_18_io_wr_instr_mem4 = io_wr_instr_mem4_18; // @[BP.scala 334:31]
  assign array_18_io_wr_instr_mem5 = io_wr_instr_mem5_18; // @[BP.scala 335:31]
  assign array_18_io_wr_instr_mem6 = io_wr_instr_mem6_18; // @[BP.scala 336:31]
  assign array_18_io_PC1_in = array_17_io_PC6_out; // @[BP.scala 338:24]
  assign array_18_io_Addr_in = array_17_io_Addr_out; // @[BP.scala 339:25]
  assign array_19_clock = clock;
  assign array_19_reset = reset;
  assign array_19_io_d_in_0_a = array_18_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_0_valid_a = array_18_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_0_b = array_18_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_0_valid_b = array_18_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_1_a = array_18_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_1_valid_a = array_18_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_1_b = array_18_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_1_valid_b = array_18_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_2_a = array_18_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_2_valid_a = array_18_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_2_b = array_18_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_2_valid_b = array_18_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_3_a = array_18_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_3_valid_a = array_18_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_3_b = array_18_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_3_valid_b = array_18_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_4_a = array_18_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_4_valid_a = array_18_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_4_b = array_18_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_4_valid_b = array_18_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_5_a = array_18_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_5_valid_a = array_18_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_5_b = array_18_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_5_valid_b = array_18_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_6_a = array_18_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_6_valid_a = array_18_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_6_b = array_18_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_6_valid_b = array_18_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_7_a = array_18_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_7_valid_a = array_18_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_7_b = array_18_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_7_valid_b = array_18_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_8_a = array_18_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_8_valid_a = array_18_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_8_b = array_18_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_8_valid_b = array_18_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_9_a = array_18_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_9_valid_a = array_18_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_9_b = array_18_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_9_valid_b = array_18_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_10_a = array_18_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_10_valid_a = array_18_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_10_b = array_18_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_10_valid_b = array_18_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_11_a = array_18_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_11_valid_a = array_18_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_11_b = array_18_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_11_valid_b = array_18_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_12_a = array_18_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_12_valid_a = array_18_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_12_b = array_18_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_12_valid_b = array_18_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_13_a = array_18_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_13_valid_a = array_18_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_13_b = array_18_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_13_valid_b = array_18_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_14_a = array_18_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_14_valid_a = array_18_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_14_b = array_18_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_14_valid_b = array_18_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_15_a = array_18_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_15_valid_a = array_18_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_15_b = array_18_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_15_valid_b = array_18_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_16_a = array_18_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_16_valid_a = array_18_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_16_b = array_18_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_16_valid_b = array_18_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_17_a = array_18_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_17_valid_a = array_18_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_17_b = array_18_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_17_valid_b = array_18_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_18_a = array_18_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_18_valid_a = array_18_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_18_b = array_18_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_18_valid_b = array_18_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_19_a = array_18_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_19_valid_a = array_18_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_19_b = array_18_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_19_valid_b = array_18_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_20_a = array_18_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_20_valid_a = array_18_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_20_b = array_18_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_20_valid_b = array_18_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_21_a = array_18_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_21_valid_a = array_18_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_21_b = array_18_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_21_valid_b = array_18_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_22_a = array_18_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_22_valid_a = array_18_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_22_b = array_18_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_22_valid_b = array_18_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_23_a = array_18_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_23_valid_a = array_18_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_23_b = array_18_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_23_valid_b = array_18_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_24_a = array_18_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_24_valid_a = array_18_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_24_b = array_18_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_24_valid_b = array_18_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_25_a = array_18_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_25_valid_a = array_18_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_25_b = array_18_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_25_valid_b = array_18_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_26_a = array_18_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_26_valid_a = array_18_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_26_b = array_18_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_26_valid_b = array_18_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_27_a = array_18_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_27_valid_a = array_18_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_27_b = array_18_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_27_valid_b = array_18_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_28_a = array_18_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_28_valid_a = array_18_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_28_b = array_18_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_28_valid_b = array_18_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_29_a = array_18_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_29_valid_a = array_18_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_29_b = array_18_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_29_valid_b = array_18_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_30_a = array_18_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_30_valid_a = array_18_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_30_b = array_18_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_30_valid_b = array_18_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_31_a = array_18_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_31_valid_a = array_18_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_19_io_d_in_31_b = array_18_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_19_io_d_in_31_valid_b = array_18_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_19_io_wr_en_mem1 = io_wr_en_mem1_19; // @[BP.scala 325:28]
  assign array_19_io_wr_en_mem2 = io_wr_en_mem2_19; // @[BP.scala 326:28]
  assign array_19_io_wr_en_mem3 = io_wr_en_mem3_19; // @[BP.scala 327:28]
  assign array_19_io_wr_en_mem4 = io_wr_en_mem4_19; // @[BP.scala 328:28]
  assign array_19_io_wr_en_mem5 = io_wr_en_mem5_19; // @[BP.scala 329:28]
  assign array_19_io_wr_en_mem6 = io_wr_en_mem6_19; // @[BP.scala 330:28]
  assign array_19_io_wr_instr_mem1 = io_wr_instr_mem1_19; // @[BP.scala 331:31]
  assign array_19_io_wr_instr_mem2 = io_wr_instr_mem2_19; // @[BP.scala 332:31]
  assign array_19_io_wr_instr_mem3 = io_wr_instr_mem3_19; // @[BP.scala 333:31]
  assign array_19_io_wr_instr_mem4 = io_wr_instr_mem4_19; // @[BP.scala 334:31]
  assign array_19_io_wr_instr_mem5 = io_wr_instr_mem5_19; // @[BP.scala 335:31]
  assign array_19_io_wr_instr_mem6 = io_wr_instr_mem6_19; // @[BP.scala 336:31]
  assign array_19_io_PC1_in = array_18_io_PC6_out; // @[BP.scala 338:24]
  assign array_19_io_Addr_in = array_18_io_Addr_out; // @[BP.scala 339:25]
  assign array_20_clock = clock;
  assign array_20_reset = reset;
  assign array_20_io_d_in_0_a = array_19_io_d_out_0_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_0_valid_a = array_19_io_d_out_0_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_0_b = array_19_io_d_out_0_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_0_valid_b = array_19_io_d_out_0_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_1_a = array_19_io_d_out_1_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_1_valid_a = array_19_io_d_out_1_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_1_b = array_19_io_d_out_1_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_1_valid_b = array_19_io_d_out_1_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_2_a = array_19_io_d_out_2_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_2_valid_a = array_19_io_d_out_2_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_2_b = array_19_io_d_out_2_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_2_valid_b = array_19_io_d_out_2_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_3_a = array_19_io_d_out_3_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_3_valid_a = array_19_io_d_out_3_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_3_b = array_19_io_d_out_3_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_3_valid_b = array_19_io_d_out_3_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_4_a = array_19_io_d_out_4_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_4_valid_a = array_19_io_d_out_4_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_4_b = array_19_io_d_out_4_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_4_valid_b = array_19_io_d_out_4_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_5_a = array_19_io_d_out_5_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_5_valid_a = array_19_io_d_out_5_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_5_b = array_19_io_d_out_5_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_5_valid_b = array_19_io_d_out_5_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_6_a = array_19_io_d_out_6_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_6_valid_a = array_19_io_d_out_6_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_6_b = array_19_io_d_out_6_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_6_valid_b = array_19_io_d_out_6_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_7_a = array_19_io_d_out_7_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_7_valid_a = array_19_io_d_out_7_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_7_b = array_19_io_d_out_7_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_7_valid_b = array_19_io_d_out_7_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_8_a = array_19_io_d_out_8_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_8_valid_a = array_19_io_d_out_8_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_8_b = array_19_io_d_out_8_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_8_valid_b = array_19_io_d_out_8_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_9_a = array_19_io_d_out_9_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_9_valid_a = array_19_io_d_out_9_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_9_b = array_19_io_d_out_9_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_9_valid_b = array_19_io_d_out_9_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_10_a = array_19_io_d_out_10_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_10_valid_a = array_19_io_d_out_10_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_10_b = array_19_io_d_out_10_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_10_valid_b = array_19_io_d_out_10_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_11_a = array_19_io_d_out_11_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_11_valid_a = array_19_io_d_out_11_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_11_b = array_19_io_d_out_11_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_11_valid_b = array_19_io_d_out_11_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_12_a = array_19_io_d_out_12_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_12_valid_a = array_19_io_d_out_12_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_12_b = array_19_io_d_out_12_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_12_valid_b = array_19_io_d_out_12_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_13_a = array_19_io_d_out_13_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_13_valid_a = array_19_io_d_out_13_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_13_b = array_19_io_d_out_13_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_13_valid_b = array_19_io_d_out_13_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_14_a = array_19_io_d_out_14_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_14_valid_a = array_19_io_d_out_14_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_14_b = array_19_io_d_out_14_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_14_valid_b = array_19_io_d_out_14_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_15_a = array_19_io_d_out_15_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_15_valid_a = array_19_io_d_out_15_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_15_b = array_19_io_d_out_15_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_15_valid_b = array_19_io_d_out_15_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_16_a = array_19_io_d_out_16_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_16_valid_a = array_19_io_d_out_16_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_16_b = array_19_io_d_out_16_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_16_valid_b = array_19_io_d_out_16_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_17_a = array_19_io_d_out_17_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_17_valid_a = array_19_io_d_out_17_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_17_b = array_19_io_d_out_17_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_17_valid_b = array_19_io_d_out_17_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_18_a = array_19_io_d_out_18_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_18_valid_a = array_19_io_d_out_18_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_18_b = array_19_io_d_out_18_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_18_valid_b = array_19_io_d_out_18_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_19_a = array_19_io_d_out_19_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_19_valid_a = array_19_io_d_out_19_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_19_b = array_19_io_d_out_19_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_19_valid_b = array_19_io_d_out_19_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_20_a = array_19_io_d_out_20_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_20_valid_a = array_19_io_d_out_20_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_20_b = array_19_io_d_out_20_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_20_valid_b = array_19_io_d_out_20_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_21_a = array_19_io_d_out_21_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_21_valid_a = array_19_io_d_out_21_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_21_b = array_19_io_d_out_21_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_21_valid_b = array_19_io_d_out_21_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_22_a = array_19_io_d_out_22_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_22_valid_a = array_19_io_d_out_22_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_22_b = array_19_io_d_out_22_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_22_valid_b = array_19_io_d_out_22_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_23_a = array_19_io_d_out_23_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_23_valid_a = array_19_io_d_out_23_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_23_b = array_19_io_d_out_23_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_23_valid_b = array_19_io_d_out_23_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_24_a = array_19_io_d_out_24_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_24_valid_a = array_19_io_d_out_24_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_24_b = array_19_io_d_out_24_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_24_valid_b = array_19_io_d_out_24_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_25_a = array_19_io_d_out_25_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_25_valid_a = array_19_io_d_out_25_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_25_b = array_19_io_d_out_25_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_25_valid_b = array_19_io_d_out_25_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_26_a = array_19_io_d_out_26_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_26_valid_a = array_19_io_d_out_26_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_26_b = array_19_io_d_out_26_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_26_valid_b = array_19_io_d_out_26_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_27_a = array_19_io_d_out_27_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_27_valid_a = array_19_io_d_out_27_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_27_b = array_19_io_d_out_27_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_27_valid_b = array_19_io_d_out_27_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_28_a = array_19_io_d_out_28_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_28_valid_a = array_19_io_d_out_28_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_28_b = array_19_io_d_out_28_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_28_valid_b = array_19_io_d_out_28_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_29_a = array_19_io_d_out_29_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_29_valid_a = array_19_io_d_out_29_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_29_b = array_19_io_d_out_29_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_29_valid_b = array_19_io_d_out_29_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_30_a = array_19_io_d_out_30_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_30_valid_a = array_19_io_d_out_30_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_30_b = array_19_io_d_out_30_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_30_valid_b = array_19_io_d_out_30_valid_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_31_a = array_19_io_d_out_31_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_31_valid_a = array_19_io_d_out_31_valid_a; // @[BP.scala 323:22]
  assign array_20_io_d_in_31_b = array_19_io_d_out_31_b; // @[BP.scala 323:22]
  assign array_20_io_d_in_31_valid_b = array_19_io_d_out_31_valid_b; // @[BP.scala 323:22]
  assign array_20_io_wr_en_mem1 = io_wr_en_mem1_20; // @[BP.scala 325:28]
  assign array_20_io_wr_en_mem2 = io_wr_en_mem2_20; // @[BP.scala 326:28]
  assign array_20_io_wr_en_mem3 = io_wr_en_mem3_20; // @[BP.scala 327:28]
  assign array_20_io_wr_en_mem4 = io_wr_en_mem4_20; // @[BP.scala 328:28]
  assign array_20_io_wr_en_mem5 = io_wr_en_mem5_20; // @[BP.scala 329:28]
  assign array_20_io_wr_en_mem6 = io_wr_en_mem6_20; // @[BP.scala 330:28]
  assign array_20_io_wr_instr_mem1 = io_wr_instr_mem1_20; // @[BP.scala 331:31]
  assign array_20_io_wr_instr_mem2 = io_wr_instr_mem2_20; // @[BP.scala 332:31]
  assign array_20_io_wr_instr_mem3 = io_wr_instr_mem3_20; // @[BP.scala 333:31]
  assign array_20_io_wr_instr_mem4 = io_wr_instr_mem4_20; // @[BP.scala 334:31]
  assign array_20_io_wr_instr_mem5 = io_wr_instr_mem5_20; // @[BP.scala 335:31]
  assign array_20_io_wr_instr_mem6 = io_wr_instr_mem6_20; // @[BP.scala 336:31]
  assign array_20_io_PC1_in = array_19_io_PC6_out; // @[BP.scala 338:24]
  assign array_20_io_Addr_in = array_19_io_Addr_out; // @[BP.scala 339:25]
  always @(posedge clock) begin
    if(inputDataBuffer_0_validBit_MPORT_en & inputDataBuffer_0_validBit_MPORT_mask) begin
      inputDataBuffer_0_validBit[inputDataBuffer_0_validBit_MPORT_addr] <= inputDataBuffer_0_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_0_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_0_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_0_data_MPORT_en & inputDataBuffer_0_data_MPORT_mask) begin
      inputDataBuffer_0_data[inputDataBuffer_0_data_MPORT_addr] <= inputDataBuffer_0_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_0_data_MPORT_3_en_pipe_0 <= io_beginRun;
    //if (io_beginRun) begin
      //inputDataBuffer_0_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    //end
    inputDataBuffer_0_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    if(inputDataBuffer_1_validBit_MPORT_en & inputDataBuffer_1_validBit_MPORT_mask) begin
      inputDataBuffer_1_validBit[inputDataBuffer_1_validBit_MPORT_addr] <= inputDataBuffer_1_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_1_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_1_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_1_data_MPORT_en & inputDataBuffer_1_data_MPORT_mask) begin
      inputDataBuffer_1_data[inputDataBuffer_1_data_MPORT_addr] <= inputDataBuffer_1_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_1_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_1_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_2_validBit_MPORT_en & inputDataBuffer_2_validBit_MPORT_mask) begin
      inputDataBuffer_2_validBit[inputDataBuffer_2_validBit_MPORT_addr] <= inputDataBuffer_2_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_2_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_2_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_2_data_MPORT_en & inputDataBuffer_2_data_MPORT_mask) begin
      inputDataBuffer_2_data[inputDataBuffer_2_data_MPORT_addr] <= inputDataBuffer_2_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_2_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_2_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_3_validBit_MPORT_en & inputDataBuffer_3_validBit_MPORT_mask) begin
      inputDataBuffer_3_validBit[inputDataBuffer_3_validBit_MPORT_addr] <= inputDataBuffer_3_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_3_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_3_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_3_data_MPORT_en & inputDataBuffer_3_data_MPORT_mask) begin
      inputDataBuffer_3_data[inputDataBuffer_3_data_MPORT_addr] <= inputDataBuffer_3_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_3_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_3_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_4_validBit_MPORT_en & inputDataBuffer_4_validBit_MPORT_mask) begin
      inputDataBuffer_4_validBit[inputDataBuffer_4_validBit_MPORT_addr] <= inputDataBuffer_4_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_4_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_4_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_4_data_MPORT_en & inputDataBuffer_4_data_MPORT_mask) begin
      inputDataBuffer_4_data[inputDataBuffer_4_data_MPORT_addr] <= inputDataBuffer_4_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_4_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_4_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_5_validBit_MPORT_en & inputDataBuffer_5_validBit_MPORT_mask) begin
      inputDataBuffer_5_validBit[inputDataBuffer_5_validBit_MPORT_addr] <= inputDataBuffer_5_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_5_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_5_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_5_data_MPORT_en & inputDataBuffer_5_data_MPORT_mask) begin
      inputDataBuffer_5_data[inputDataBuffer_5_data_MPORT_addr] <= inputDataBuffer_5_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_5_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_5_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_6_validBit_MPORT_en & inputDataBuffer_6_validBit_MPORT_mask) begin
      inputDataBuffer_6_validBit[inputDataBuffer_6_validBit_MPORT_addr] <= inputDataBuffer_6_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_6_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_6_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_6_data_MPORT_en & inputDataBuffer_6_data_MPORT_mask) begin
      inputDataBuffer_6_data[inputDataBuffer_6_data_MPORT_addr] <= inputDataBuffer_6_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_6_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_6_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_7_validBit_MPORT_en & inputDataBuffer_7_validBit_MPORT_mask) begin
      inputDataBuffer_7_validBit[inputDataBuffer_7_validBit_MPORT_addr] <= inputDataBuffer_7_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_7_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_7_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_7_data_MPORT_en & inputDataBuffer_7_data_MPORT_mask) begin
      inputDataBuffer_7_data[inputDataBuffer_7_data_MPORT_addr] <= inputDataBuffer_7_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_7_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_7_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_8_validBit_MPORT_en & inputDataBuffer_8_validBit_MPORT_mask) begin
      inputDataBuffer_8_validBit[inputDataBuffer_8_validBit_MPORT_addr] <= inputDataBuffer_8_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_8_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_8_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_8_data_MPORT_en & inputDataBuffer_8_data_MPORT_mask) begin
      inputDataBuffer_8_data[inputDataBuffer_8_data_MPORT_addr] <= inputDataBuffer_8_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_8_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_8_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_9_validBit_MPORT_en & inputDataBuffer_9_validBit_MPORT_mask) begin
      inputDataBuffer_9_validBit[inputDataBuffer_9_validBit_MPORT_addr] <= inputDataBuffer_9_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_9_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_9_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_9_data_MPORT_en & inputDataBuffer_9_data_MPORT_mask) begin
      inputDataBuffer_9_data[inputDataBuffer_9_data_MPORT_addr] <= inputDataBuffer_9_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_9_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_9_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_10_validBit_MPORT_en & inputDataBuffer_10_validBit_MPORT_mask) begin
      inputDataBuffer_10_validBit[inputDataBuffer_10_validBit_MPORT_addr] <= inputDataBuffer_10_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_10_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_10_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_10_data_MPORT_en & inputDataBuffer_10_data_MPORT_mask) begin
      inputDataBuffer_10_data[inputDataBuffer_10_data_MPORT_addr] <= inputDataBuffer_10_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_10_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_10_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_11_validBit_MPORT_en & inputDataBuffer_11_validBit_MPORT_mask) begin
      inputDataBuffer_11_validBit[inputDataBuffer_11_validBit_MPORT_addr] <= inputDataBuffer_11_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_11_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_11_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_11_data_MPORT_en & inputDataBuffer_11_data_MPORT_mask) begin
      inputDataBuffer_11_data[inputDataBuffer_11_data_MPORT_addr] <= inputDataBuffer_11_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_11_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_11_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_12_validBit_MPORT_en & inputDataBuffer_12_validBit_MPORT_mask) begin
      inputDataBuffer_12_validBit[inputDataBuffer_12_validBit_MPORT_addr] <= inputDataBuffer_12_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_12_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_12_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_12_data_MPORT_en & inputDataBuffer_12_data_MPORT_mask) begin
      inputDataBuffer_12_data[inputDataBuffer_12_data_MPORT_addr] <= inputDataBuffer_12_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_12_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_12_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_13_validBit_MPORT_en & inputDataBuffer_13_validBit_MPORT_mask) begin
      inputDataBuffer_13_validBit[inputDataBuffer_13_validBit_MPORT_addr] <= inputDataBuffer_13_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_13_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_13_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_13_data_MPORT_en & inputDataBuffer_13_data_MPORT_mask) begin
      inputDataBuffer_13_data[inputDataBuffer_13_data_MPORT_addr] <= inputDataBuffer_13_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_13_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_13_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_14_validBit_MPORT_en & inputDataBuffer_14_validBit_MPORT_mask) begin
      inputDataBuffer_14_validBit[inputDataBuffer_14_validBit_MPORT_addr] <= inputDataBuffer_14_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_14_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_14_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_14_data_MPORT_en & inputDataBuffer_14_data_MPORT_mask) begin
      inputDataBuffer_14_data[inputDataBuffer_14_data_MPORT_addr] <= inputDataBuffer_14_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_14_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_14_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_15_validBit_MPORT_en & inputDataBuffer_15_validBit_MPORT_mask) begin
      inputDataBuffer_15_validBit[inputDataBuffer_15_validBit_MPORT_addr] <= inputDataBuffer_15_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_15_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_15_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_15_data_MPORT_en & inputDataBuffer_15_data_MPORT_mask) begin
      inputDataBuffer_15_data[inputDataBuffer_15_data_MPORT_addr] <= inputDataBuffer_15_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_15_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_15_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_16_validBit_MPORT_en & inputDataBuffer_16_validBit_MPORT_mask) begin
      inputDataBuffer_16_validBit[inputDataBuffer_16_validBit_MPORT_addr] <= inputDataBuffer_16_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_16_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_16_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_16_data_MPORT_en & inputDataBuffer_16_data_MPORT_mask) begin
      inputDataBuffer_16_data[inputDataBuffer_16_data_MPORT_addr] <= inputDataBuffer_16_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_16_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_16_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_17_validBit_MPORT_en & inputDataBuffer_17_validBit_MPORT_mask) begin
      inputDataBuffer_17_validBit[inputDataBuffer_17_validBit_MPORT_addr] <= inputDataBuffer_17_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_17_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_17_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_17_data_MPORT_en & inputDataBuffer_17_data_MPORT_mask) begin
      inputDataBuffer_17_data[inputDataBuffer_17_data_MPORT_addr] <= inputDataBuffer_17_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_17_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_17_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_18_validBit_MPORT_en & inputDataBuffer_18_validBit_MPORT_mask) begin
      inputDataBuffer_18_validBit[inputDataBuffer_18_validBit_MPORT_addr] <= inputDataBuffer_18_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_18_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_18_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_18_data_MPORT_en & inputDataBuffer_18_data_MPORT_mask) begin
      inputDataBuffer_18_data[inputDataBuffer_18_data_MPORT_addr] <= inputDataBuffer_18_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_18_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_18_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_19_validBit_MPORT_en & inputDataBuffer_19_validBit_MPORT_mask) begin
      inputDataBuffer_19_validBit[inputDataBuffer_19_validBit_MPORT_addr] <= inputDataBuffer_19_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_19_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_19_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_19_data_MPORT_en & inputDataBuffer_19_data_MPORT_mask) begin
      inputDataBuffer_19_data[inputDataBuffer_19_data_MPORT_addr] <= inputDataBuffer_19_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_19_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_19_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_20_validBit_MPORT_en & inputDataBuffer_20_validBit_MPORT_mask) begin
      inputDataBuffer_20_validBit[inputDataBuffer_20_validBit_MPORT_addr] <= inputDataBuffer_20_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_20_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_20_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_20_data_MPORT_en & inputDataBuffer_20_data_MPORT_mask) begin
      inputDataBuffer_20_data[inputDataBuffer_20_data_MPORT_addr] <= inputDataBuffer_20_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_20_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_20_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_21_validBit_MPORT_en & inputDataBuffer_21_validBit_MPORT_mask) begin
      inputDataBuffer_21_validBit[inputDataBuffer_21_validBit_MPORT_addr] <= inputDataBuffer_21_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_21_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_21_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_21_data_MPORT_en & inputDataBuffer_21_data_MPORT_mask) begin
      inputDataBuffer_21_data[inputDataBuffer_21_data_MPORT_addr] <= inputDataBuffer_21_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_21_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_21_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_22_validBit_MPORT_en & inputDataBuffer_22_validBit_MPORT_mask) begin
      inputDataBuffer_22_validBit[inputDataBuffer_22_validBit_MPORT_addr] <= inputDataBuffer_22_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_22_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_22_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_22_data_MPORT_en & inputDataBuffer_22_data_MPORT_mask) begin
      inputDataBuffer_22_data[inputDataBuffer_22_data_MPORT_addr] <= inputDataBuffer_22_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_22_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_22_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_23_validBit_MPORT_en & inputDataBuffer_23_validBit_MPORT_mask) begin
      inputDataBuffer_23_validBit[inputDataBuffer_23_validBit_MPORT_addr] <= inputDataBuffer_23_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_23_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_23_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_23_data_MPORT_en & inputDataBuffer_23_data_MPORT_mask) begin
      inputDataBuffer_23_data[inputDataBuffer_23_data_MPORT_addr] <= inputDataBuffer_23_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_23_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_23_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_24_validBit_MPORT_en & inputDataBuffer_24_validBit_MPORT_mask) begin
      inputDataBuffer_24_validBit[inputDataBuffer_24_validBit_MPORT_addr] <= inputDataBuffer_24_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_24_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_24_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_24_data_MPORT_en & inputDataBuffer_24_data_MPORT_mask) begin
      inputDataBuffer_24_data[inputDataBuffer_24_data_MPORT_addr] <= inputDataBuffer_24_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_24_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_24_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_25_validBit_MPORT_en & inputDataBuffer_25_validBit_MPORT_mask) begin
      inputDataBuffer_25_validBit[inputDataBuffer_25_validBit_MPORT_addr] <= inputDataBuffer_25_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_25_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_25_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_25_data_MPORT_en & inputDataBuffer_25_data_MPORT_mask) begin
      inputDataBuffer_25_data[inputDataBuffer_25_data_MPORT_addr] <= inputDataBuffer_25_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_25_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_25_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_26_validBit_MPORT_en & inputDataBuffer_26_validBit_MPORT_mask) begin
      inputDataBuffer_26_validBit[inputDataBuffer_26_validBit_MPORT_addr] <= inputDataBuffer_26_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_26_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_26_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_26_data_MPORT_en & inputDataBuffer_26_data_MPORT_mask) begin
      inputDataBuffer_26_data[inputDataBuffer_26_data_MPORT_addr] <= inputDataBuffer_26_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_26_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_26_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_27_validBit_MPORT_en & inputDataBuffer_27_validBit_MPORT_mask) begin
      inputDataBuffer_27_validBit[inputDataBuffer_27_validBit_MPORT_addr] <= inputDataBuffer_27_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_27_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_27_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_27_data_MPORT_en & inputDataBuffer_27_data_MPORT_mask) begin
      inputDataBuffer_27_data[inputDataBuffer_27_data_MPORT_addr] <= inputDataBuffer_27_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_27_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_27_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_28_validBit_MPORT_en & inputDataBuffer_28_validBit_MPORT_mask) begin
      inputDataBuffer_28_validBit[inputDataBuffer_28_validBit_MPORT_addr] <= inputDataBuffer_28_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_28_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_28_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_28_data_MPORT_en & inputDataBuffer_28_data_MPORT_mask) begin
      inputDataBuffer_28_data[inputDataBuffer_28_data_MPORT_addr] <= inputDataBuffer_28_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_28_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_28_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_29_validBit_MPORT_en & inputDataBuffer_29_validBit_MPORT_mask) begin
      inputDataBuffer_29_validBit[inputDataBuffer_29_validBit_MPORT_addr] <= inputDataBuffer_29_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_29_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_29_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_29_data_MPORT_en & inputDataBuffer_29_data_MPORT_mask) begin
      inputDataBuffer_29_data[inputDataBuffer_29_data_MPORT_addr] <= inputDataBuffer_29_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_29_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_29_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_30_validBit_MPORT_en & inputDataBuffer_30_validBit_MPORT_mask) begin
      inputDataBuffer_30_validBit[inputDataBuffer_30_validBit_MPORT_addr] <= inputDataBuffer_30_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_30_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_30_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_30_data_MPORT_en & inputDataBuffer_30_data_MPORT_mask) begin
      inputDataBuffer_30_data[inputDataBuffer_30_data_MPORT_addr] <= inputDataBuffer_30_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_30_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_30_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_31_validBit_MPORT_en & inputDataBuffer_31_validBit_MPORT_mask) begin
      inputDataBuffer_31_validBit[inputDataBuffer_31_validBit_MPORT_addr] <= inputDataBuffer_31_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_31_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_31_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_31_data_MPORT_en & inputDataBuffer_31_data_MPORT_mask) begin
      inputDataBuffer_31_data[inputDataBuffer_31_data_MPORT_addr] <= inputDataBuffer_31_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_31_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_31_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_32_validBit_MPORT_en & inputDataBuffer_32_validBit_MPORT_mask) begin
      inputDataBuffer_32_validBit[inputDataBuffer_32_validBit_MPORT_addr] <= inputDataBuffer_32_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_32_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_32_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_32_data_MPORT_en & inputDataBuffer_32_data_MPORT_mask) begin
      inputDataBuffer_32_data[inputDataBuffer_32_data_MPORT_addr] <= inputDataBuffer_32_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_32_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_32_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_33_validBit_MPORT_en & inputDataBuffer_33_validBit_MPORT_mask) begin
      inputDataBuffer_33_validBit[inputDataBuffer_33_validBit_MPORT_addr] <= inputDataBuffer_33_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_33_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_33_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_33_data_MPORT_en & inputDataBuffer_33_data_MPORT_mask) begin
      inputDataBuffer_33_data[inputDataBuffer_33_data_MPORT_addr] <= inputDataBuffer_33_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_33_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_33_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_34_validBit_MPORT_en & inputDataBuffer_34_validBit_MPORT_mask) begin
      inputDataBuffer_34_validBit[inputDataBuffer_34_validBit_MPORT_addr] <= inputDataBuffer_34_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_34_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_34_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_34_data_MPORT_en & inputDataBuffer_34_data_MPORT_mask) begin
      inputDataBuffer_34_data[inputDataBuffer_34_data_MPORT_addr] <= inputDataBuffer_34_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_34_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_34_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_35_validBit_MPORT_en & inputDataBuffer_35_validBit_MPORT_mask) begin
      inputDataBuffer_35_validBit[inputDataBuffer_35_validBit_MPORT_addr] <= inputDataBuffer_35_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_35_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_35_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_35_data_MPORT_en & inputDataBuffer_35_data_MPORT_mask) begin
      inputDataBuffer_35_data[inputDataBuffer_35_data_MPORT_addr] <= inputDataBuffer_35_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_35_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_35_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_36_validBit_MPORT_en & inputDataBuffer_36_validBit_MPORT_mask) begin
      inputDataBuffer_36_validBit[inputDataBuffer_36_validBit_MPORT_addr] <= inputDataBuffer_36_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_36_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_36_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_36_data_MPORT_en & inputDataBuffer_36_data_MPORT_mask) begin
      inputDataBuffer_36_data[inputDataBuffer_36_data_MPORT_addr] <= inputDataBuffer_36_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_36_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_36_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_37_validBit_MPORT_en & inputDataBuffer_37_validBit_MPORT_mask) begin
      inputDataBuffer_37_validBit[inputDataBuffer_37_validBit_MPORT_addr] <= inputDataBuffer_37_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_37_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_37_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_37_data_MPORT_en & inputDataBuffer_37_data_MPORT_mask) begin
      inputDataBuffer_37_data[inputDataBuffer_37_data_MPORT_addr] <= inputDataBuffer_37_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_37_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_37_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_38_validBit_MPORT_en & inputDataBuffer_38_validBit_MPORT_mask) begin
      inputDataBuffer_38_validBit[inputDataBuffer_38_validBit_MPORT_addr] <= inputDataBuffer_38_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_38_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_38_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_38_data_MPORT_en & inputDataBuffer_38_data_MPORT_mask) begin
      inputDataBuffer_38_data[inputDataBuffer_38_data_MPORT_addr] <= inputDataBuffer_38_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_38_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_38_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_39_validBit_MPORT_en & inputDataBuffer_39_validBit_MPORT_mask) begin
      inputDataBuffer_39_validBit[inputDataBuffer_39_validBit_MPORT_addr] <= inputDataBuffer_39_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_39_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_39_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_39_data_MPORT_en & inputDataBuffer_39_data_MPORT_mask) begin
      inputDataBuffer_39_data[inputDataBuffer_39_data_MPORT_addr] <= inputDataBuffer_39_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_39_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_39_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_40_validBit_MPORT_en & inputDataBuffer_40_validBit_MPORT_mask) begin
      inputDataBuffer_40_validBit[inputDataBuffer_40_validBit_MPORT_addr] <= inputDataBuffer_40_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_40_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_40_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_40_data_MPORT_en & inputDataBuffer_40_data_MPORT_mask) begin
      inputDataBuffer_40_data[inputDataBuffer_40_data_MPORT_addr] <= inputDataBuffer_40_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_40_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_40_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_41_validBit_MPORT_en & inputDataBuffer_41_validBit_MPORT_mask) begin
      inputDataBuffer_41_validBit[inputDataBuffer_41_validBit_MPORT_addr] <= inputDataBuffer_41_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_41_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_41_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_41_data_MPORT_en & inputDataBuffer_41_data_MPORT_mask) begin
      inputDataBuffer_41_data[inputDataBuffer_41_data_MPORT_addr] <= inputDataBuffer_41_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_41_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_41_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_42_validBit_MPORT_en & inputDataBuffer_42_validBit_MPORT_mask) begin
      inputDataBuffer_42_validBit[inputDataBuffer_42_validBit_MPORT_addr] <= inputDataBuffer_42_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_42_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_42_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_42_data_MPORT_en & inputDataBuffer_42_data_MPORT_mask) begin
      inputDataBuffer_42_data[inputDataBuffer_42_data_MPORT_addr] <= inputDataBuffer_42_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_42_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_42_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_43_validBit_MPORT_en & inputDataBuffer_43_validBit_MPORT_mask) begin
      inputDataBuffer_43_validBit[inputDataBuffer_43_validBit_MPORT_addr] <= inputDataBuffer_43_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_43_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_43_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_43_data_MPORT_en & inputDataBuffer_43_data_MPORT_mask) begin
      inputDataBuffer_43_data[inputDataBuffer_43_data_MPORT_addr] <= inputDataBuffer_43_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_43_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_43_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_44_validBit_MPORT_en & inputDataBuffer_44_validBit_MPORT_mask) begin
      inputDataBuffer_44_validBit[inputDataBuffer_44_validBit_MPORT_addr] <= inputDataBuffer_44_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_44_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_44_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_44_data_MPORT_en & inputDataBuffer_44_data_MPORT_mask) begin
      inputDataBuffer_44_data[inputDataBuffer_44_data_MPORT_addr] <= inputDataBuffer_44_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_44_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_44_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_45_validBit_MPORT_en & inputDataBuffer_45_validBit_MPORT_mask) begin
      inputDataBuffer_45_validBit[inputDataBuffer_45_validBit_MPORT_addr] <= inputDataBuffer_45_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_45_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_45_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_45_data_MPORT_en & inputDataBuffer_45_data_MPORT_mask) begin
      inputDataBuffer_45_data[inputDataBuffer_45_data_MPORT_addr] <= inputDataBuffer_45_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_45_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_45_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_46_validBit_MPORT_en & inputDataBuffer_46_validBit_MPORT_mask) begin
      inputDataBuffer_46_validBit[inputDataBuffer_46_validBit_MPORT_addr] <= inputDataBuffer_46_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_46_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_46_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_46_data_MPORT_en & inputDataBuffer_46_data_MPORT_mask) begin
      inputDataBuffer_46_data[inputDataBuffer_46_data_MPORT_addr] <= inputDataBuffer_46_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_46_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_46_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_47_validBit_MPORT_en & inputDataBuffer_47_validBit_MPORT_mask) begin
      inputDataBuffer_47_validBit[inputDataBuffer_47_validBit_MPORT_addr] <= inputDataBuffer_47_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_47_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_47_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_47_data_MPORT_en & inputDataBuffer_47_data_MPORT_mask) begin
      inputDataBuffer_47_data[inputDataBuffer_47_data_MPORT_addr] <= inputDataBuffer_47_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_47_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_47_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_48_validBit_MPORT_en & inputDataBuffer_48_validBit_MPORT_mask) begin
      inputDataBuffer_48_validBit[inputDataBuffer_48_validBit_MPORT_addr] <= inputDataBuffer_48_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_48_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_48_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_48_data_MPORT_en & inputDataBuffer_48_data_MPORT_mask) begin
      inputDataBuffer_48_data[inputDataBuffer_48_data_MPORT_addr] <= inputDataBuffer_48_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_48_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_48_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_49_validBit_MPORT_en & inputDataBuffer_49_validBit_MPORT_mask) begin
      inputDataBuffer_49_validBit[inputDataBuffer_49_validBit_MPORT_addr] <= inputDataBuffer_49_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_49_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_49_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_49_data_MPORT_en & inputDataBuffer_49_data_MPORT_mask) begin
      inputDataBuffer_49_data[inputDataBuffer_49_data_MPORT_addr] <= inputDataBuffer_49_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_49_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_49_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_50_validBit_MPORT_en & inputDataBuffer_50_validBit_MPORT_mask) begin
      inputDataBuffer_50_validBit[inputDataBuffer_50_validBit_MPORT_addr] <= inputDataBuffer_50_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_50_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_50_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_50_data_MPORT_en & inputDataBuffer_50_data_MPORT_mask) begin
      inputDataBuffer_50_data[inputDataBuffer_50_data_MPORT_addr] <= inputDataBuffer_50_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_50_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_50_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_51_validBit_MPORT_en & inputDataBuffer_51_validBit_MPORT_mask) begin
      inputDataBuffer_51_validBit[inputDataBuffer_51_validBit_MPORT_addr] <= inputDataBuffer_51_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_51_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_51_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_51_data_MPORT_en & inputDataBuffer_51_data_MPORT_mask) begin
      inputDataBuffer_51_data[inputDataBuffer_51_data_MPORT_addr] <= inputDataBuffer_51_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_51_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_51_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_52_validBit_MPORT_en & inputDataBuffer_52_validBit_MPORT_mask) begin
      inputDataBuffer_52_validBit[inputDataBuffer_52_validBit_MPORT_addr] <= inputDataBuffer_52_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_52_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_52_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_52_data_MPORT_en & inputDataBuffer_52_data_MPORT_mask) begin
      inputDataBuffer_52_data[inputDataBuffer_52_data_MPORT_addr] <= inputDataBuffer_52_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_52_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_52_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_53_validBit_MPORT_en & inputDataBuffer_53_validBit_MPORT_mask) begin
      inputDataBuffer_53_validBit[inputDataBuffer_53_validBit_MPORT_addr] <= inputDataBuffer_53_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_53_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_53_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_53_data_MPORT_en & inputDataBuffer_53_data_MPORT_mask) begin
      inputDataBuffer_53_data[inputDataBuffer_53_data_MPORT_addr] <= inputDataBuffer_53_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_53_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_53_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_54_validBit_MPORT_en & inputDataBuffer_54_validBit_MPORT_mask) begin
      inputDataBuffer_54_validBit[inputDataBuffer_54_validBit_MPORT_addr] <= inputDataBuffer_54_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_54_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_54_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_54_data_MPORT_en & inputDataBuffer_54_data_MPORT_mask) begin
      inputDataBuffer_54_data[inputDataBuffer_54_data_MPORT_addr] <= inputDataBuffer_54_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_54_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_54_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_55_validBit_MPORT_en & inputDataBuffer_55_validBit_MPORT_mask) begin
      inputDataBuffer_55_validBit[inputDataBuffer_55_validBit_MPORT_addr] <= inputDataBuffer_55_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_55_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_55_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_55_data_MPORT_en & inputDataBuffer_55_data_MPORT_mask) begin
      inputDataBuffer_55_data[inputDataBuffer_55_data_MPORT_addr] <= inputDataBuffer_55_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_55_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_55_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_56_validBit_MPORT_en & inputDataBuffer_56_validBit_MPORT_mask) begin
      inputDataBuffer_56_validBit[inputDataBuffer_56_validBit_MPORT_addr] <= inputDataBuffer_56_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_56_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_56_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_56_data_MPORT_en & inputDataBuffer_56_data_MPORT_mask) begin
      inputDataBuffer_56_data[inputDataBuffer_56_data_MPORT_addr] <= inputDataBuffer_56_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_56_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_56_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_57_validBit_MPORT_en & inputDataBuffer_57_validBit_MPORT_mask) begin
      inputDataBuffer_57_validBit[inputDataBuffer_57_validBit_MPORT_addr] <= inputDataBuffer_57_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_57_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_57_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_57_data_MPORT_en & inputDataBuffer_57_data_MPORT_mask) begin
      inputDataBuffer_57_data[inputDataBuffer_57_data_MPORT_addr] <= inputDataBuffer_57_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_57_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_57_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_58_validBit_MPORT_en & inputDataBuffer_58_validBit_MPORT_mask) begin
      inputDataBuffer_58_validBit[inputDataBuffer_58_validBit_MPORT_addr] <= inputDataBuffer_58_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_58_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_58_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_58_data_MPORT_en & inputDataBuffer_58_data_MPORT_mask) begin
      inputDataBuffer_58_data[inputDataBuffer_58_data_MPORT_addr] <= inputDataBuffer_58_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_58_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_58_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_59_validBit_MPORT_en & inputDataBuffer_59_validBit_MPORT_mask) begin
      inputDataBuffer_59_validBit[inputDataBuffer_59_validBit_MPORT_addr] <= inputDataBuffer_59_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_59_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_59_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_59_data_MPORT_en & inputDataBuffer_59_data_MPORT_mask) begin
      inputDataBuffer_59_data[inputDataBuffer_59_data_MPORT_addr] <= inputDataBuffer_59_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_59_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_59_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_60_validBit_MPORT_en & inputDataBuffer_60_validBit_MPORT_mask) begin
      inputDataBuffer_60_validBit[inputDataBuffer_60_validBit_MPORT_addr] <= inputDataBuffer_60_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_60_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_60_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_60_data_MPORT_en & inputDataBuffer_60_data_MPORT_mask) begin
      inputDataBuffer_60_data[inputDataBuffer_60_data_MPORT_addr] <= inputDataBuffer_60_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_60_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_60_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_61_validBit_MPORT_en & inputDataBuffer_61_validBit_MPORT_mask) begin
      inputDataBuffer_61_validBit[inputDataBuffer_61_validBit_MPORT_addr] <= inputDataBuffer_61_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_61_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_61_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_61_data_MPORT_en & inputDataBuffer_61_data_MPORT_mask) begin
      inputDataBuffer_61_data[inputDataBuffer_61_data_MPORT_addr] <= inputDataBuffer_61_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_61_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_61_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_62_validBit_MPORT_en & inputDataBuffer_62_validBit_MPORT_mask) begin
      inputDataBuffer_62_validBit[inputDataBuffer_62_validBit_MPORT_addr] <= inputDataBuffer_62_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_62_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_62_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_62_data_MPORT_en & inputDataBuffer_62_data_MPORT_mask) begin
      inputDataBuffer_62_data[inputDataBuffer_62_data_MPORT_addr] <= inputDataBuffer_62_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_62_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_62_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_63_validBit_MPORT_en & inputDataBuffer_63_validBit_MPORT_mask) begin
      inputDataBuffer_63_validBit[inputDataBuffer_63_validBit_MPORT_addr] <= inputDataBuffer_63_validBit_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_63_validBit_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_63_validBit_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(inputDataBuffer_63_data_MPORT_en & inputDataBuffer_63_data_MPORT_mask) begin
      inputDataBuffer_63_data[inputDataBuffer_63_data_MPORT_addr] <= inputDataBuffer_63_data_MPORT_data; // @[BP.scala 42:36]
    end
    inputDataBuffer_63_data_MPORT_3_en_pipe_0 <= io_beginRun;
    if (io_beginRun) begin
      inputDataBuffer_63_data_MPORT_3_addr_pipe_0 <= rd_Addr_inBuf;
    end
    if(outputDataBuffer_0_validBit_MPORT_4_en & outputDataBuffer_0_validBit_MPORT_4_mask) begin
      outputDataBuffer_0_validBit[outputDataBuffer_0_validBit_MPORT_4_addr] <= outputDataBuffer_0_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_0_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_0_data_MPORT_4_en & outputDataBuffer_0_data_MPORT_4_mask) begin
      outputDataBuffer_0_data[outputDataBuffer_0_data_MPORT_4_addr] <= outputDataBuffer_0_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_0_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_1_validBit_MPORT_4_en & outputDataBuffer_1_validBit_MPORT_4_mask) begin
      outputDataBuffer_1_validBit[outputDataBuffer_1_validBit_MPORT_4_addr] <= outputDataBuffer_1_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_1_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_1_data_MPORT_4_en & outputDataBuffer_1_data_MPORT_4_mask) begin
      outputDataBuffer_1_data[outputDataBuffer_1_data_MPORT_4_addr] <= outputDataBuffer_1_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_1_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_2_validBit_MPORT_4_en & outputDataBuffer_2_validBit_MPORT_4_mask) begin
      outputDataBuffer_2_validBit[outputDataBuffer_2_validBit_MPORT_4_addr] <= outputDataBuffer_2_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_2_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_2_data_MPORT_4_en & outputDataBuffer_2_data_MPORT_4_mask) begin
      outputDataBuffer_2_data[outputDataBuffer_2_data_MPORT_4_addr] <= outputDataBuffer_2_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_2_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_3_validBit_MPORT_4_en & outputDataBuffer_3_validBit_MPORT_4_mask) begin
      outputDataBuffer_3_validBit[outputDataBuffer_3_validBit_MPORT_4_addr] <= outputDataBuffer_3_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_3_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_3_data_MPORT_4_en & outputDataBuffer_3_data_MPORT_4_mask) begin
      outputDataBuffer_3_data[outputDataBuffer_3_data_MPORT_4_addr] <= outputDataBuffer_3_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_3_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_4_validBit_MPORT_4_en & outputDataBuffer_4_validBit_MPORT_4_mask) begin
      outputDataBuffer_4_validBit[outputDataBuffer_4_validBit_MPORT_4_addr] <= outputDataBuffer_4_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_4_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_4_data_MPORT_4_en & outputDataBuffer_4_data_MPORT_4_mask) begin
      outputDataBuffer_4_data[outputDataBuffer_4_data_MPORT_4_addr] <= outputDataBuffer_4_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_4_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_5_validBit_MPORT_4_en & outputDataBuffer_5_validBit_MPORT_4_mask) begin
      outputDataBuffer_5_validBit[outputDataBuffer_5_validBit_MPORT_4_addr] <= outputDataBuffer_5_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_5_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_5_data_MPORT_4_en & outputDataBuffer_5_data_MPORT_4_mask) begin
      outputDataBuffer_5_data[outputDataBuffer_5_data_MPORT_4_addr] <= outputDataBuffer_5_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_5_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_6_validBit_MPORT_4_en & outputDataBuffer_6_validBit_MPORT_4_mask) begin
      outputDataBuffer_6_validBit[outputDataBuffer_6_validBit_MPORT_4_addr] <= outputDataBuffer_6_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_6_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_6_data_MPORT_4_en & outputDataBuffer_6_data_MPORT_4_mask) begin
      outputDataBuffer_6_data[outputDataBuffer_6_data_MPORT_4_addr] <= outputDataBuffer_6_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_6_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_7_validBit_MPORT_4_en & outputDataBuffer_7_validBit_MPORT_4_mask) begin
      outputDataBuffer_7_validBit[outputDataBuffer_7_validBit_MPORT_4_addr] <= outputDataBuffer_7_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_7_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_7_data_MPORT_4_en & outputDataBuffer_7_data_MPORT_4_mask) begin
      outputDataBuffer_7_data[outputDataBuffer_7_data_MPORT_4_addr] <= outputDataBuffer_7_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_7_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_8_validBit_MPORT_4_en & outputDataBuffer_8_validBit_MPORT_4_mask) begin
      outputDataBuffer_8_validBit[outputDataBuffer_8_validBit_MPORT_4_addr] <= outputDataBuffer_8_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_8_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_8_data_MPORT_4_en & outputDataBuffer_8_data_MPORT_4_mask) begin
      outputDataBuffer_8_data[outputDataBuffer_8_data_MPORT_4_addr] <= outputDataBuffer_8_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_8_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_9_validBit_MPORT_4_en & outputDataBuffer_9_validBit_MPORT_4_mask) begin
      outputDataBuffer_9_validBit[outputDataBuffer_9_validBit_MPORT_4_addr] <= outputDataBuffer_9_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_9_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_9_data_MPORT_4_en & outputDataBuffer_9_data_MPORT_4_mask) begin
      outputDataBuffer_9_data[outputDataBuffer_9_data_MPORT_4_addr] <= outputDataBuffer_9_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_9_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_10_validBit_MPORT_4_en & outputDataBuffer_10_validBit_MPORT_4_mask) begin
      outputDataBuffer_10_validBit[outputDataBuffer_10_validBit_MPORT_4_addr] <=
        outputDataBuffer_10_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_10_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_10_data_MPORT_4_en & outputDataBuffer_10_data_MPORT_4_mask) begin
      outputDataBuffer_10_data[outputDataBuffer_10_data_MPORT_4_addr] <= outputDataBuffer_10_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_10_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_11_validBit_MPORT_4_en & outputDataBuffer_11_validBit_MPORT_4_mask) begin
      outputDataBuffer_11_validBit[outputDataBuffer_11_validBit_MPORT_4_addr] <=
        outputDataBuffer_11_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_11_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_11_data_MPORT_4_en & outputDataBuffer_11_data_MPORT_4_mask) begin
      outputDataBuffer_11_data[outputDataBuffer_11_data_MPORT_4_addr] <= outputDataBuffer_11_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_11_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_12_validBit_MPORT_4_en & outputDataBuffer_12_validBit_MPORT_4_mask) begin
      outputDataBuffer_12_validBit[outputDataBuffer_12_validBit_MPORT_4_addr] <=
        outputDataBuffer_12_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_12_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_12_data_MPORT_4_en & outputDataBuffer_12_data_MPORT_4_mask) begin
      outputDataBuffer_12_data[outputDataBuffer_12_data_MPORT_4_addr] <= outputDataBuffer_12_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_12_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_13_validBit_MPORT_4_en & outputDataBuffer_13_validBit_MPORT_4_mask) begin
      outputDataBuffer_13_validBit[outputDataBuffer_13_validBit_MPORT_4_addr] <=
        outputDataBuffer_13_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_13_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_13_data_MPORT_4_en & outputDataBuffer_13_data_MPORT_4_mask) begin
      outputDataBuffer_13_data[outputDataBuffer_13_data_MPORT_4_addr] <= outputDataBuffer_13_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_13_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_14_validBit_MPORT_4_en & outputDataBuffer_14_validBit_MPORT_4_mask) begin
      outputDataBuffer_14_validBit[outputDataBuffer_14_validBit_MPORT_4_addr] <=
        outputDataBuffer_14_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_14_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_14_data_MPORT_4_en & outputDataBuffer_14_data_MPORT_4_mask) begin
      outputDataBuffer_14_data[outputDataBuffer_14_data_MPORT_4_addr] <= outputDataBuffer_14_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_14_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_15_validBit_MPORT_4_en & outputDataBuffer_15_validBit_MPORT_4_mask) begin
      outputDataBuffer_15_validBit[outputDataBuffer_15_validBit_MPORT_4_addr] <=
        outputDataBuffer_15_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_15_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_15_data_MPORT_4_en & outputDataBuffer_15_data_MPORT_4_mask) begin
      outputDataBuffer_15_data[outputDataBuffer_15_data_MPORT_4_addr] <= outputDataBuffer_15_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_15_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_16_validBit_MPORT_4_en & outputDataBuffer_16_validBit_MPORT_4_mask) begin
      outputDataBuffer_16_validBit[outputDataBuffer_16_validBit_MPORT_4_addr] <=
        outputDataBuffer_16_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_16_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_16_data_MPORT_4_en & outputDataBuffer_16_data_MPORT_4_mask) begin
      outputDataBuffer_16_data[outputDataBuffer_16_data_MPORT_4_addr] <= outputDataBuffer_16_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_16_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_17_validBit_MPORT_4_en & outputDataBuffer_17_validBit_MPORT_4_mask) begin
      outputDataBuffer_17_validBit[outputDataBuffer_17_validBit_MPORT_4_addr] <=
        outputDataBuffer_17_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_17_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_17_data_MPORT_4_en & outputDataBuffer_17_data_MPORT_4_mask) begin
      outputDataBuffer_17_data[outputDataBuffer_17_data_MPORT_4_addr] <= outputDataBuffer_17_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_17_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_18_validBit_MPORT_4_en & outputDataBuffer_18_validBit_MPORT_4_mask) begin
      outputDataBuffer_18_validBit[outputDataBuffer_18_validBit_MPORT_4_addr] <=
        outputDataBuffer_18_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_18_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_18_data_MPORT_4_en & outputDataBuffer_18_data_MPORT_4_mask) begin
      outputDataBuffer_18_data[outputDataBuffer_18_data_MPORT_4_addr] <= outputDataBuffer_18_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_18_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_19_validBit_MPORT_4_en & outputDataBuffer_19_validBit_MPORT_4_mask) begin
      outputDataBuffer_19_validBit[outputDataBuffer_19_validBit_MPORT_4_addr] <=
        outputDataBuffer_19_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_19_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_19_data_MPORT_4_en & outputDataBuffer_19_data_MPORT_4_mask) begin
      outputDataBuffer_19_data[outputDataBuffer_19_data_MPORT_4_addr] <= outputDataBuffer_19_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_19_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_20_validBit_MPORT_4_en & outputDataBuffer_20_validBit_MPORT_4_mask) begin
      outputDataBuffer_20_validBit[outputDataBuffer_20_validBit_MPORT_4_addr] <=
        outputDataBuffer_20_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_20_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_20_data_MPORT_4_en & outputDataBuffer_20_data_MPORT_4_mask) begin
      outputDataBuffer_20_data[outputDataBuffer_20_data_MPORT_4_addr] <= outputDataBuffer_20_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_20_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_21_validBit_MPORT_4_en & outputDataBuffer_21_validBit_MPORT_4_mask) begin
      outputDataBuffer_21_validBit[outputDataBuffer_21_validBit_MPORT_4_addr] <=
        outputDataBuffer_21_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_21_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_21_data_MPORT_4_en & outputDataBuffer_21_data_MPORT_4_mask) begin
      outputDataBuffer_21_data[outputDataBuffer_21_data_MPORT_4_addr] <= outputDataBuffer_21_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_21_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_22_validBit_MPORT_4_en & outputDataBuffer_22_validBit_MPORT_4_mask) begin
      outputDataBuffer_22_validBit[outputDataBuffer_22_validBit_MPORT_4_addr] <=
        outputDataBuffer_22_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_22_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_22_data_MPORT_4_en & outputDataBuffer_22_data_MPORT_4_mask) begin
      outputDataBuffer_22_data[outputDataBuffer_22_data_MPORT_4_addr] <= outputDataBuffer_22_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_22_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_23_validBit_MPORT_4_en & outputDataBuffer_23_validBit_MPORT_4_mask) begin
      outputDataBuffer_23_validBit[outputDataBuffer_23_validBit_MPORT_4_addr] <=
        outputDataBuffer_23_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_23_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_23_data_MPORT_4_en & outputDataBuffer_23_data_MPORT_4_mask) begin
      outputDataBuffer_23_data[outputDataBuffer_23_data_MPORT_4_addr] <= outputDataBuffer_23_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_23_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_24_validBit_MPORT_4_en & outputDataBuffer_24_validBit_MPORT_4_mask) begin
      outputDataBuffer_24_validBit[outputDataBuffer_24_validBit_MPORT_4_addr] <=
        outputDataBuffer_24_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_24_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_24_data_MPORT_4_en & outputDataBuffer_24_data_MPORT_4_mask) begin
      outputDataBuffer_24_data[outputDataBuffer_24_data_MPORT_4_addr] <= outputDataBuffer_24_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_24_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_25_validBit_MPORT_4_en & outputDataBuffer_25_validBit_MPORT_4_mask) begin
      outputDataBuffer_25_validBit[outputDataBuffer_25_validBit_MPORT_4_addr] <=
        outputDataBuffer_25_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_25_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_25_data_MPORT_4_en & outputDataBuffer_25_data_MPORT_4_mask) begin
      outputDataBuffer_25_data[outputDataBuffer_25_data_MPORT_4_addr] <= outputDataBuffer_25_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_25_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_26_validBit_MPORT_4_en & outputDataBuffer_26_validBit_MPORT_4_mask) begin
      outputDataBuffer_26_validBit[outputDataBuffer_26_validBit_MPORT_4_addr] <=
        outputDataBuffer_26_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_26_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_26_data_MPORT_4_en & outputDataBuffer_26_data_MPORT_4_mask) begin
      outputDataBuffer_26_data[outputDataBuffer_26_data_MPORT_4_addr] <= outputDataBuffer_26_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_26_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_27_validBit_MPORT_4_en & outputDataBuffer_27_validBit_MPORT_4_mask) begin
      outputDataBuffer_27_validBit[outputDataBuffer_27_validBit_MPORT_4_addr] <=
        outputDataBuffer_27_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_27_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_27_data_MPORT_4_en & outputDataBuffer_27_data_MPORT_4_mask) begin
      outputDataBuffer_27_data[outputDataBuffer_27_data_MPORT_4_addr] <= outputDataBuffer_27_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_27_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_28_validBit_MPORT_4_en & outputDataBuffer_28_validBit_MPORT_4_mask) begin
      outputDataBuffer_28_validBit[outputDataBuffer_28_validBit_MPORT_4_addr] <=
        outputDataBuffer_28_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_28_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_28_data_MPORT_4_en & outputDataBuffer_28_data_MPORT_4_mask) begin
      outputDataBuffer_28_data[outputDataBuffer_28_data_MPORT_4_addr] <= outputDataBuffer_28_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_28_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_29_validBit_MPORT_4_en & outputDataBuffer_29_validBit_MPORT_4_mask) begin
      outputDataBuffer_29_validBit[outputDataBuffer_29_validBit_MPORT_4_addr] <=
        outputDataBuffer_29_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_29_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_29_data_MPORT_4_en & outputDataBuffer_29_data_MPORT_4_mask) begin
      outputDataBuffer_29_data[outputDataBuffer_29_data_MPORT_4_addr] <= outputDataBuffer_29_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_29_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_30_validBit_MPORT_4_en & outputDataBuffer_30_validBit_MPORT_4_mask) begin
      outputDataBuffer_30_validBit[outputDataBuffer_30_validBit_MPORT_4_addr] <=
        outputDataBuffer_30_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_30_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_30_data_MPORT_4_en & outputDataBuffer_30_data_MPORT_4_mask) begin
      outputDataBuffer_30_data[outputDataBuffer_30_data_MPORT_4_addr] <= outputDataBuffer_30_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_30_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_31_validBit_MPORT_4_en & outputDataBuffer_31_validBit_MPORT_4_mask) begin
      outputDataBuffer_31_validBit[outputDataBuffer_31_validBit_MPORT_4_addr] <=
        outputDataBuffer_31_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_31_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_31_data_MPORT_4_en & outputDataBuffer_31_data_MPORT_4_mask) begin
      outputDataBuffer_31_data[outputDataBuffer_31_data_MPORT_4_addr] <= outputDataBuffer_31_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_31_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_32_validBit_MPORT_4_en & outputDataBuffer_32_validBit_MPORT_4_mask) begin
      outputDataBuffer_32_validBit[outputDataBuffer_32_validBit_MPORT_4_addr] <=
        outputDataBuffer_32_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_32_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_32_data_MPORT_4_en & outputDataBuffer_32_data_MPORT_4_mask) begin
      outputDataBuffer_32_data[outputDataBuffer_32_data_MPORT_4_addr] <= outputDataBuffer_32_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_32_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_33_validBit_MPORT_4_en & outputDataBuffer_33_validBit_MPORT_4_mask) begin
      outputDataBuffer_33_validBit[outputDataBuffer_33_validBit_MPORT_4_addr] <=
        outputDataBuffer_33_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_33_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_33_data_MPORT_4_en & outputDataBuffer_33_data_MPORT_4_mask) begin
      outputDataBuffer_33_data[outputDataBuffer_33_data_MPORT_4_addr] <= outputDataBuffer_33_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_33_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_34_validBit_MPORT_4_en & outputDataBuffer_34_validBit_MPORT_4_mask) begin
      outputDataBuffer_34_validBit[outputDataBuffer_34_validBit_MPORT_4_addr] <=
        outputDataBuffer_34_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_34_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_34_data_MPORT_4_en & outputDataBuffer_34_data_MPORT_4_mask) begin
      outputDataBuffer_34_data[outputDataBuffer_34_data_MPORT_4_addr] <= outputDataBuffer_34_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_34_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_35_validBit_MPORT_4_en & outputDataBuffer_35_validBit_MPORT_4_mask) begin
      outputDataBuffer_35_validBit[outputDataBuffer_35_validBit_MPORT_4_addr] <=
        outputDataBuffer_35_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_35_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_35_data_MPORT_4_en & outputDataBuffer_35_data_MPORT_4_mask) begin
      outputDataBuffer_35_data[outputDataBuffer_35_data_MPORT_4_addr] <= outputDataBuffer_35_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_35_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_36_validBit_MPORT_4_en & outputDataBuffer_36_validBit_MPORT_4_mask) begin
      outputDataBuffer_36_validBit[outputDataBuffer_36_validBit_MPORT_4_addr] <=
        outputDataBuffer_36_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_36_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_36_data_MPORT_4_en & outputDataBuffer_36_data_MPORT_4_mask) begin
      outputDataBuffer_36_data[outputDataBuffer_36_data_MPORT_4_addr] <= outputDataBuffer_36_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_36_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_37_validBit_MPORT_4_en & outputDataBuffer_37_validBit_MPORT_4_mask) begin
      outputDataBuffer_37_validBit[outputDataBuffer_37_validBit_MPORT_4_addr] <=
        outputDataBuffer_37_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_37_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_37_data_MPORT_4_en & outputDataBuffer_37_data_MPORT_4_mask) begin
      outputDataBuffer_37_data[outputDataBuffer_37_data_MPORT_4_addr] <= outputDataBuffer_37_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_37_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_38_validBit_MPORT_4_en & outputDataBuffer_38_validBit_MPORT_4_mask) begin
      outputDataBuffer_38_validBit[outputDataBuffer_38_validBit_MPORT_4_addr] <=
        outputDataBuffer_38_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_38_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_38_data_MPORT_4_en & outputDataBuffer_38_data_MPORT_4_mask) begin
      outputDataBuffer_38_data[outputDataBuffer_38_data_MPORT_4_addr] <= outputDataBuffer_38_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_38_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_39_validBit_MPORT_4_en & outputDataBuffer_39_validBit_MPORT_4_mask) begin
      outputDataBuffer_39_validBit[outputDataBuffer_39_validBit_MPORT_4_addr] <=
        outputDataBuffer_39_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_39_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_39_data_MPORT_4_en & outputDataBuffer_39_data_MPORT_4_mask) begin
      outputDataBuffer_39_data[outputDataBuffer_39_data_MPORT_4_addr] <= outputDataBuffer_39_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_39_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_40_validBit_MPORT_4_en & outputDataBuffer_40_validBit_MPORT_4_mask) begin
      outputDataBuffer_40_validBit[outputDataBuffer_40_validBit_MPORT_4_addr] <=
        outputDataBuffer_40_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_40_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_40_data_MPORT_4_en & outputDataBuffer_40_data_MPORT_4_mask) begin
      outputDataBuffer_40_data[outputDataBuffer_40_data_MPORT_4_addr] <= outputDataBuffer_40_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_40_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_41_validBit_MPORT_4_en & outputDataBuffer_41_validBit_MPORT_4_mask) begin
      outputDataBuffer_41_validBit[outputDataBuffer_41_validBit_MPORT_4_addr] <=
        outputDataBuffer_41_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_41_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_41_data_MPORT_4_en & outputDataBuffer_41_data_MPORT_4_mask) begin
      outputDataBuffer_41_data[outputDataBuffer_41_data_MPORT_4_addr] <= outputDataBuffer_41_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_41_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_42_validBit_MPORT_4_en & outputDataBuffer_42_validBit_MPORT_4_mask) begin
      outputDataBuffer_42_validBit[outputDataBuffer_42_validBit_MPORT_4_addr] <=
        outputDataBuffer_42_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_42_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_42_data_MPORT_4_en & outputDataBuffer_42_data_MPORT_4_mask) begin
      outputDataBuffer_42_data[outputDataBuffer_42_data_MPORT_4_addr] <= outputDataBuffer_42_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_42_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_43_validBit_MPORT_4_en & outputDataBuffer_43_validBit_MPORT_4_mask) begin
      outputDataBuffer_43_validBit[outputDataBuffer_43_validBit_MPORT_4_addr] <=
        outputDataBuffer_43_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_43_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_43_data_MPORT_4_en & outputDataBuffer_43_data_MPORT_4_mask) begin
      outputDataBuffer_43_data[outputDataBuffer_43_data_MPORT_4_addr] <= outputDataBuffer_43_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_43_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_44_validBit_MPORT_4_en & outputDataBuffer_44_validBit_MPORT_4_mask) begin
      outputDataBuffer_44_validBit[outputDataBuffer_44_validBit_MPORT_4_addr] <=
        outputDataBuffer_44_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_44_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_44_data_MPORT_4_en & outputDataBuffer_44_data_MPORT_4_mask) begin
      outputDataBuffer_44_data[outputDataBuffer_44_data_MPORT_4_addr] <= outputDataBuffer_44_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_44_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_45_validBit_MPORT_4_en & outputDataBuffer_45_validBit_MPORT_4_mask) begin
      outputDataBuffer_45_validBit[outputDataBuffer_45_validBit_MPORT_4_addr] <=
        outputDataBuffer_45_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_45_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_45_data_MPORT_4_en & outputDataBuffer_45_data_MPORT_4_mask) begin
      outputDataBuffer_45_data[outputDataBuffer_45_data_MPORT_4_addr] <= outputDataBuffer_45_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_45_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_46_validBit_MPORT_4_en & outputDataBuffer_46_validBit_MPORT_4_mask) begin
      outputDataBuffer_46_validBit[outputDataBuffer_46_validBit_MPORT_4_addr] <=
        outputDataBuffer_46_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_46_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_46_data_MPORT_4_en & outputDataBuffer_46_data_MPORT_4_mask) begin
      outputDataBuffer_46_data[outputDataBuffer_46_data_MPORT_4_addr] <= outputDataBuffer_46_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_46_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_47_validBit_MPORT_4_en & outputDataBuffer_47_validBit_MPORT_4_mask) begin
      outputDataBuffer_47_validBit[outputDataBuffer_47_validBit_MPORT_4_addr] <=
        outputDataBuffer_47_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_47_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_47_data_MPORT_4_en & outputDataBuffer_47_data_MPORT_4_mask) begin
      outputDataBuffer_47_data[outputDataBuffer_47_data_MPORT_4_addr] <= outputDataBuffer_47_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_47_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_48_validBit_MPORT_4_en & outputDataBuffer_48_validBit_MPORT_4_mask) begin
      outputDataBuffer_48_validBit[outputDataBuffer_48_validBit_MPORT_4_addr] <=
        outputDataBuffer_48_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_48_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_48_data_MPORT_4_en & outputDataBuffer_48_data_MPORT_4_mask) begin
      outputDataBuffer_48_data[outputDataBuffer_48_data_MPORT_4_addr] <= outputDataBuffer_48_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_48_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_49_validBit_MPORT_4_en & outputDataBuffer_49_validBit_MPORT_4_mask) begin
      outputDataBuffer_49_validBit[outputDataBuffer_49_validBit_MPORT_4_addr] <=
        outputDataBuffer_49_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_49_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_49_data_MPORT_4_en & outputDataBuffer_49_data_MPORT_4_mask) begin
      outputDataBuffer_49_data[outputDataBuffer_49_data_MPORT_4_addr] <= outputDataBuffer_49_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_49_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_50_validBit_MPORT_4_en & outputDataBuffer_50_validBit_MPORT_4_mask) begin
      outputDataBuffer_50_validBit[outputDataBuffer_50_validBit_MPORT_4_addr] <=
        outputDataBuffer_50_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_50_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_50_data_MPORT_4_en & outputDataBuffer_50_data_MPORT_4_mask) begin
      outputDataBuffer_50_data[outputDataBuffer_50_data_MPORT_4_addr] <= outputDataBuffer_50_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_50_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_51_validBit_MPORT_4_en & outputDataBuffer_51_validBit_MPORT_4_mask) begin
      outputDataBuffer_51_validBit[outputDataBuffer_51_validBit_MPORT_4_addr] <=
        outputDataBuffer_51_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_51_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_51_data_MPORT_4_en & outputDataBuffer_51_data_MPORT_4_mask) begin
      outputDataBuffer_51_data[outputDataBuffer_51_data_MPORT_4_addr] <= outputDataBuffer_51_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_51_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_52_validBit_MPORT_4_en & outputDataBuffer_52_validBit_MPORT_4_mask) begin
      outputDataBuffer_52_validBit[outputDataBuffer_52_validBit_MPORT_4_addr] <=
        outputDataBuffer_52_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_52_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_52_data_MPORT_4_en & outputDataBuffer_52_data_MPORT_4_mask) begin
      outputDataBuffer_52_data[outputDataBuffer_52_data_MPORT_4_addr] <= outputDataBuffer_52_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_52_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_53_validBit_MPORT_4_en & outputDataBuffer_53_validBit_MPORT_4_mask) begin
      outputDataBuffer_53_validBit[outputDataBuffer_53_validBit_MPORT_4_addr] <=
        outputDataBuffer_53_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_53_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_53_data_MPORT_4_en & outputDataBuffer_53_data_MPORT_4_mask) begin
      outputDataBuffer_53_data[outputDataBuffer_53_data_MPORT_4_addr] <= outputDataBuffer_53_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_53_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_54_validBit_MPORT_4_en & outputDataBuffer_54_validBit_MPORT_4_mask) begin
      outputDataBuffer_54_validBit[outputDataBuffer_54_validBit_MPORT_4_addr] <=
        outputDataBuffer_54_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_54_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_54_data_MPORT_4_en & outputDataBuffer_54_data_MPORT_4_mask) begin
      outputDataBuffer_54_data[outputDataBuffer_54_data_MPORT_4_addr] <= outputDataBuffer_54_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_54_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_55_validBit_MPORT_4_en & outputDataBuffer_55_validBit_MPORT_4_mask) begin
      outputDataBuffer_55_validBit[outputDataBuffer_55_validBit_MPORT_4_addr] <=
        outputDataBuffer_55_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_55_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_55_data_MPORT_4_en & outputDataBuffer_55_data_MPORT_4_mask) begin
      outputDataBuffer_55_data[outputDataBuffer_55_data_MPORT_4_addr] <= outputDataBuffer_55_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_55_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_56_validBit_MPORT_4_en & outputDataBuffer_56_validBit_MPORT_4_mask) begin
      outputDataBuffer_56_validBit[outputDataBuffer_56_validBit_MPORT_4_addr] <=
        outputDataBuffer_56_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_56_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_56_data_MPORT_4_en & outputDataBuffer_56_data_MPORT_4_mask) begin
      outputDataBuffer_56_data[outputDataBuffer_56_data_MPORT_4_addr] <= outputDataBuffer_56_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_56_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_57_validBit_MPORT_4_en & outputDataBuffer_57_validBit_MPORT_4_mask) begin
      outputDataBuffer_57_validBit[outputDataBuffer_57_validBit_MPORT_4_addr] <=
        outputDataBuffer_57_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_57_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_57_data_MPORT_4_en & outputDataBuffer_57_data_MPORT_4_mask) begin
      outputDataBuffer_57_data[outputDataBuffer_57_data_MPORT_4_addr] <= outputDataBuffer_57_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_57_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_58_validBit_MPORT_4_en & outputDataBuffer_58_validBit_MPORT_4_mask) begin
      outputDataBuffer_58_validBit[outputDataBuffer_58_validBit_MPORT_4_addr] <=
        outputDataBuffer_58_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_58_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_58_data_MPORT_4_en & outputDataBuffer_58_data_MPORT_4_mask) begin
      outputDataBuffer_58_data[outputDataBuffer_58_data_MPORT_4_addr] <= outputDataBuffer_58_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_58_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_59_validBit_MPORT_4_en & outputDataBuffer_59_validBit_MPORT_4_mask) begin
      outputDataBuffer_59_validBit[outputDataBuffer_59_validBit_MPORT_4_addr] <=
        outputDataBuffer_59_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_59_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_59_data_MPORT_4_en & outputDataBuffer_59_data_MPORT_4_mask) begin
      outputDataBuffer_59_data[outputDataBuffer_59_data_MPORT_4_addr] <= outputDataBuffer_59_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_59_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_60_validBit_MPORT_4_en & outputDataBuffer_60_validBit_MPORT_4_mask) begin
      outputDataBuffer_60_validBit[outputDataBuffer_60_validBit_MPORT_4_addr] <=
        outputDataBuffer_60_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_60_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_60_data_MPORT_4_en & outputDataBuffer_60_data_MPORT_4_mask) begin
      outputDataBuffer_60_data[outputDataBuffer_60_data_MPORT_4_addr] <= outputDataBuffer_60_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_60_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_61_validBit_MPORT_4_en & outputDataBuffer_61_validBit_MPORT_4_mask) begin
      outputDataBuffer_61_validBit[outputDataBuffer_61_validBit_MPORT_4_addr] <=
        outputDataBuffer_61_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_61_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_61_data_MPORT_4_en & outputDataBuffer_61_data_MPORT_4_mask) begin
      outputDataBuffer_61_data[outputDataBuffer_61_data_MPORT_4_addr] <= outputDataBuffer_61_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_61_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_62_validBit_MPORT_4_en & outputDataBuffer_62_validBit_MPORT_4_mask) begin
      outputDataBuffer_62_validBit[outputDataBuffer_62_validBit_MPORT_4_addr] <=
        outputDataBuffer_62_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_62_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_62_data_MPORT_4_en & outputDataBuffer_62_data_MPORT_4_mask) begin
      outputDataBuffer_62_data[outputDataBuffer_62_data_MPORT_4_addr] <= outputDataBuffer_62_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_62_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_63_validBit_MPORT_4_en & outputDataBuffer_63_validBit_MPORT_4_mask) begin
      outputDataBuffer_63_validBit[outputDataBuffer_63_validBit_MPORT_4_addr] <=
        outputDataBuffer_63_validBit_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_63_validBit_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if(outputDataBuffer_63_data_MPORT_4_en & outputDataBuffer_63_data_MPORT_4_mask) begin
      outputDataBuffer_63_data[outputDataBuffer_63_data_MPORT_4_addr] <= outputDataBuffer_63_data_MPORT_4_data; // @[BP.scala 47:37]
    end
    outputDataBuffer_63_data_MPORT_2_addr_pipe_0 <= io_rd_Addr_outBuf;
    if (reset) begin // @[BP.scala 50:30]
      wr_Addr_inBuf <= 8'h0; // @[BP.scala 50:30]
    end else if (io_wr_Addr_inBuf_en) begin // @[BP.scala 58:28]
      wr_Addr_inBuf <= _wr_Addr_inBuf_T_1; // @[BP.scala 61:19]
    end
    if (reset) begin // @[BP.scala 91:30]
      rd_Addr_inBuf <= 8'h0; // @[BP.scala 91:30]
    end else if (io_beginRun) begin // @[BP.scala 100:20]
      rd_Addr_inBuf <= _rd_Addr_inBuf_T_1; // @[BP.scala 101:19]
    end
    rd_D_inBuf_0_validBit <= inputDataBuffer_0_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_0_data <= inputDataBuffer_0_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_1_validBit <= inputDataBuffer_1_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_1_data <= inputDataBuffer_1_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_2_validBit <= inputDataBuffer_2_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_2_data <= inputDataBuffer_2_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_3_validBit <= inputDataBuffer_3_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_3_data <= inputDataBuffer_3_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_4_validBit <= inputDataBuffer_4_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_4_data <= inputDataBuffer_4_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_5_validBit <= inputDataBuffer_5_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_5_data <= inputDataBuffer_5_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_6_validBit <= inputDataBuffer_6_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_6_data <= inputDataBuffer_6_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_7_validBit <= inputDataBuffer_7_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_7_data <= inputDataBuffer_7_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_8_validBit <= inputDataBuffer_8_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_8_data <= inputDataBuffer_8_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_9_validBit <= inputDataBuffer_9_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_9_data <= inputDataBuffer_9_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_10_validBit <= inputDataBuffer_10_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_10_data <= inputDataBuffer_10_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_11_validBit <= inputDataBuffer_11_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_11_data <= inputDataBuffer_11_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_12_validBit <= inputDataBuffer_12_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_12_data <= inputDataBuffer_12_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_13_validBit <= inputDataBuffer_13_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_13_data <= inputDataBuffer_13_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_14_validBit <= inputDataBuffer_14_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_14_data <= inputDataBuffer_14_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_15_validBit <= inputDataBuffer_15_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_15_data <= inputDataBuffer_15_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_16_validBit <= inputDataBuffer_16_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_16_data <= inputDataBuffer_16_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_17_validBit <= inputDataBuffer_17_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_17_data <= inputDataBuffer_17_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_18_validBit <= inputDataBuffer_18_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_18_data <= inputDataBuffer_18_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_19_validBit <= inputDataBuffer_19_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_19_data <= inputDataBuffer_19_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_20_validBit <= inputDataBuffer_20_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_20_data <= inputDataBuffer_20_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_21_validBit <= inputDataBuffer_21_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_21_data <= inputDataBuffer_21_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_22_validBit <= inputDataBuffer_22_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_22_data <= inputDataBuffer_22_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_23_validBit <= inputDataBuffer_23_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_23_data <= inputDataBuffer_23_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_24_validBit <= inputDataBuffer_24_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_24_data <= inputDataBuffer_24_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_25_validBit <= inputDataBuffer_25_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_25_data <= inputDataBuffer_25_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_26_validBit <= inputDataBuffer_26_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_26_data <= inputDataBuffer_26_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_27_validBit <= inputDataBuffer_27_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_27_data <= inputDataBuffer_27_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_28_validBit <= inputDataBuffer_28_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_28_data <= inputDataBuffer_28_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_29_validBit <= inputDataBuffer_29_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_29_data <= inputDataBuffer_29_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_30_validBit <= inputDataBuffer_30_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_30_data <= inputDataBuffer_30_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_31_validBit <= inputDataBuffer_31_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_31_data <= inputDataBuffer_31_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_32_validBit <= inputDataBuffer_32_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_32_data <= inputDataBuffer_32_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_33_validBit <= inputDataBuffer_33_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_33_data <= inputDataBuffer_33_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_34_validBit <= inputDataBuffer_34_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_34_data <= inputDataBuffer_34_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_35_validBit <= inputDataBuffer_35_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_35_data <= inputDataBuffer_35_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_36_validBit <= inputDataBuffer_36_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_36_data <= inputDataBuffer_36_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_37_validBit <= inputDataBuffer_37_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_37_data <= inputDataBuffer_37_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_38_validBit <= inputDataBuffer_38_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_38_data <= inputDataBuffer_38_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_39_validBit <= inputDataBuffer_39_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_39_data <= inputDataBuffer_39_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_40_validBit <= inputDataBuffer_40_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_40_data <= inputDataBuffer_40_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_41_validBit <= inputDataBuffer_41_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_41_data <= inputDataBuffer_41_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_42_validBit <= inputDataBuffer_42_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_42_data <= inputDataBuffer_42_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_43_validBit <= inputDataBuffer_43_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_43_data <= inputDataBuffer_43_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_44_validBit <= inputDataBuffer_44_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_44_data <= inputDataBuffer_44_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_45_validBit <= inputDataBuffer_45_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_45_data <= inputDataBuffer_45_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_46_validBit <= inputDataBuffer_46_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_46_data <= inputDataBuffer_46_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_47_validBit <= inputDataBuffer_47_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_47_data <= inputDataBuffer_47_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_48_validBit <= inputDataBuffer_48_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_48_data <= inputDataBuffer_48_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_49_validBit <= inputDataBuffer_49_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_49_data <= inputDataBuffer_49_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_50_validBit <= inputDataBuffer_50_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_50_data <= inputDataBuffer_50_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_51_validBit <= inputDataBuffer_51_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_51_data <= inputDataBuffer_51_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_52_validBit <= inputDataBuffer_52_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_52_data <= inputDataBuffer_52_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_53_validBit <= inputDataBuffer_53_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_53_data <= inputDataBuffer_53_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_54_validBit <= inputDataBuffer_54_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_54_data <= inputDataBuffer_54_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_55_validBit <= inputDataBuffer_55_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_55_data <= inputDataBuffer_55_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_56_validBit <= inputDataBuffer_56_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_56_data <= inputDataBuffer_56_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_57_validBit <= inputDataBuffer_57_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_57_data <= inputDataBuffer_57_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_58_validBit <= inputDataBuffer_58_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_58_data <= inputDataBuffer_58_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_59_validBit <= inputDataBuffer_59_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_59_data <= inputDataBuffer_59_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_60_validBit <= inputDataBuffer_60_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_60_data <= inputDataBuffer_60_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_61_validBit <= inputDataBuffer_61_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_61_data <= inputDataBuffer_61_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_62_validBit <= inputDataBuffer_62_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_62_data <= inputDataBuffer_62_data_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_63_validBit <= inputDataBuffer_63_validBit_MPORT_3_data; // @[BP.scala 98:14]
    rd_D_inBuf_63_data <= inputDataBuffer_63_data_MPORT_3_data; // @[BP.scala 98:14]
    if (reset) begin // @[BP.scala 114:31]
      wr_Addr_outBuf <= 8'h0; // @[BP.scala 114:31]
    end else begin
      wr_Addr_outBuf <= Addr_out; // @[BP.scala 122:18]
    end
    wr_D_outBuf_0_validBit <= array_20_io_d_out_0_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_0_data <= array_20_io_d_out_0_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_1_validBit <= array_20_io_d_out_0_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_1_data <= array_20_io_d_out_0_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_2_validBit <= array_20_io_d_out_1_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_2_data <= array_20_io_d_out_1_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_3_validBit <= array_20_io_d_out_1_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_3_data <= array_20_io_d_out_1_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_4_validBit <= array_20_io_d_out_2_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_4_data <= array_20_io_d_out_2_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_5_validBit <= array_20_io_d_out_2_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_5_data <= array_20_io_d_out_2_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_6_validBit <= array_20_io_d_out_3_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_6_data <= array_20_io_d_out_3_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_7_validBit <= array_20_io_d_out_3_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_7_data <= array_20_io_d_out_3_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_8_validBit <= array_20_io_d_out_4_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_8_data <= array_20_io_d_out_4_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_9_validBit <= array_20_io_d_out_4_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_9_data <= array_20_io_d_out_4_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_10_validBit <= array_20_io_d_out_5_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_10_data <= array_20_io_d_out_5_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_11_validBit <= array_20_io_d_out_5_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_11_data <= array_20_io_d_out_5_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_12_validBit <= array_20_io_d_out_6_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_12_data <= array_20_io_d_out_6_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_13_validBit <= array_20_io_d_out_6_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_13_data <= array_20_io_d_out_6_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_14_validBit <= array_20_io_d_out_7_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_14_data <= array_20_io_d_out_7_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_15_validBit <= array_20_io_d_out_7_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_15_data <= array_20_io_d_out_7_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_16_validBit <= array_20_io_d_out_8_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_16_data <= array_20_io_d_out_8_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_17_validBit <= array_20_io_d_out_8_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_17_data <= array_20_io_d_out_8_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_18_validBit <= array_20_io_d_out_9_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_18_data <= array_20_io_d_out_9_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_19_validBit <= array_20_io_d_out_9_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_19_data <= array_20_io_d_out_9_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_20_validBit <= array_20_io_d_out_10_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_20_data <= array_20_io_d_out_10_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_21_validBit <= array_20_io_d_out_10_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_21_data <= array_20_io_d_out_10_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_22_validBit <= array_20_io_d_out_11_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_22_data <= array_20_io_d_out_11_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_23_validBit <= array_20_io_d_out_11_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_23_data <= array_20_io_d_out_11_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_24_validBit <= array_20_io_d_out_12_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_24_data <= array_20_io_d_out_12_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_25_validBit <= array_20_io_d_out_12_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_25_data <= array_20_io_d_out_12_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_26_validBit <= array_20_io_d_out_13_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_26_data <= array_20_io_d_out_13_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_27_validBit <= array_20_io_d_out_13_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_27_data <= array_20_io_d_out_13_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_28_validBit <= array_20_io_d_out_14_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_28_data <= array_20_io_d_out_14_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_29_validBit <= array_20_io_d_out_14_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_29_data <= array_20_io_d_out_14_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_30_validBit <= array_20_io_d_out_15_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_30_data <= array_20_io_d_out_15_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_31_validBit <= array_20_io_d_out_15_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_31_data <= array_20_io_d_out_15_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_32_validBit <= array_20_io_d_out_16_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_32_data <= array_20_io_d_out_16_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_33_validBit <= array_20_io_d_out_16_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_33_data <= array_20_io_d_out_16_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_34_validBit <= array_20_io_d_out_17_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_34_data <= array_20_io_d_out_17_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_35_validBit <= array_20_io_d_out_17_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_35_data <= array_20_io_d_out_17_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_36_validBit <= array_20_io_d_out_18_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_36_data <= array_20_io_d_out_18_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_37_validBit <= array_20_io_d_out_18_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_37_data <= array_20_io_d_out_18_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_38_validBit <= array_20_io_d_out_19_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_38_data <= array_20_io_d_out_19_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_39_validBit <= array_20_io_d_out_19_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_39_data <= array_20_io_d_out_19_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_40_validBit <= array_20_io_d_out_20_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_40_data <= array_20_io_d_out_20_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_41_validBit <= array_20_io_d_out_20_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_41_data <= array_20_io_d_out_20_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_42_validBit <= array_20_io_d_out_21_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_42_data <= array_20_io_d_out_21_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_43_validBit <= array_20_io_d_out_21_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_43_data <= array_20_io_d_out_21_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_44_validBit <= array_20_io_d_out_22_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_44_data <= array_20_io_d_out_22_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_45_validBit <= array_20_io_d_out_22_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_45_data <= array_20_io_d_out_22_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_46_validBit <= array_20_io_d_out_23_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_46_data <= array_20_io_d_out_23_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_47_validBit <= array_20_io_d_out_23_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_47_data <= array_20_io_d_out_23_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_48_validBit <= array_20_io_d_out_24_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_48_data <= array_20_io_d_out_24_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_49_validBit <= array_20_io_d_out_24_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_49_data <= array_20_io_d_out_24_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_50_validBit <= array_20_io_d_out_25_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_50_data <= array_20_io_d_out_25_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_51_validBit <= array_20_io_d_out_25_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_51_data <= array_20_io_d_out_25_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_52_validBit <= array_20_io_d_out_26_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_52_data <= array_20_io_d_out_26_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_53_validBit <= array_20_io_d_out_26_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_53_data <= array_20_io_d_out_26_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_54_validBit <= array_20_io_d_out_27_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_54_data <= array_20_io_d_out_27_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_55_validBit <= array_20_io_d_out_27_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_55_data <= array_20_io_d_out_27_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_56_validBit <= array_20_io_d_out_28_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_56_data <= array_20_io_d_out_28_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_57_validBit <= array_20_io_d_out_28_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_57_data <= array_20_io_d_out_28_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_58_validBit <= array_20_io_d_out_29_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_58_data <= array_20_io_d_out_29_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_59_validBit <= array_20_io_d_out_29_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_59_data <= array_20_io_d_out_29_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_60_validBit <= array_20_io_d_out_30_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_60_data <= array_20_io_d_out_30_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_61_validBit <= array_20_io_d_out_30_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_61_data <= array_20_io_d_out_30_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_62_validBit <= array_20_io_d_out_31_valid_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_62_data <= array_20_io_d_out_31_a; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_63_validBit <= array_20_io_d_out_31_valid_b; // @[BP.scala 230:19 BP.scala 342:9]
    wr_D_outBuf_63_data <= array_20_io_d_out_31_b; // @[BP.scala 230:19 BP.scala 342:9]
    if (reset) begin // @[BP.scala 287:24]
      PCBegin <= 8'h0; // @[BP.scala 287:24]
    end else if (io_beginRun) begin // @[BP.scala 294:21]
      PCBegin <= _PCBegin_T_1; // @[BP.scala 295:13]
    end
    if (reset) begin // @[BP.scala 288:26]
      AddrBegin <= 8'h0; // @[BP.scala 288:26]
    end else if (io_beginRun) begin // @[BP.scala 298:21]
      AddrBegin <= _AddrBegin_T_1; // @[BP.scala 299:15]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_0_validBit[initvar] = _RAND_0[0:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_0_data[initvar] = _RAND_3[3:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_1_validBit[initvar] = _RAND_6[0:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_1_data[initvar] = _RAND_9[3:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_2_validBit[initvar] = _RAND_12[0:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_2_data[initvar] = _RAND_15[3:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_3_validBit[initvar] = _RAND_18[0:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_3_data[initvar] = _RAND_21[3:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_4_validBit[initvar] = _RAND_24[0:0];
  _RAND_27 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_4_data[initvar] = _RAND_27[3:0];
  _RAND_30 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_5_validBit[initvar] = _RAND_30[0:0];
  _RAND_33 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_5_data[initvar] = _RAND_33[3:0];
  _RAND_36 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_6_validBit[initvar] = _RAND_36[0:0];
  _RAND_39 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_6_data[initvar] = _RAND_39[3:0];
  _RAND_42 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_7_validBit[initvar] = _RAND_42[0:0];
  _RAND_45 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_7_data[initvar] = _RAND_45[3:0];
  _RAND_48 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_8_validBit[initvar] = _RAND_48[0:0];
  _RAND_51 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_8_data[initvar] = _RAND_51[3:0];
  _RAND_54 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_9_validBit[initvar] = _RAND_54[0:0];
  _RAND_57 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_9_data[initvar] = _RAND_57[3:0];
  _RAND_60 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_10_validBit[initvar] = _RAND_60[0:0];
  _RAND_63 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_10_data[initvar] = _RAND_63[3:0];
  _RAND_66 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_11_validBit[initvar] = _RAND_66[0:0];
  _RAND_69 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_11_data[initvar] = _RAND_69[3:0];
  _RAND_72 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_12_validBit[initvar] = _RAND_72[0:0];
  _RAND_75 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_12_data[initvar] = _RAND_75[3:0];
  _RAND_78 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_13_validBit[initvar] = _RAND_78[0:0];
  _RAND_81 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_13_data[initvar] = _RAND_81[3:0];
  _RAND_84 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_14_validBit[initvar] = _RAND_84[0:0];
  _RAND_87 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_14_data[initvar] = _RAND_87[3:0];
  _RAND_90 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_15_validBit[initvar] = _RAND_90[0:0];
  _RAND_93 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_15_data[initvar] = _RAND_93[3:0];
  _RAND_96 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_16_validBit[initvar] = _RAND_96[0:0];
  _RAND_99 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_16_data[initvar] = _RAND_99[3:0];
  _RAND_102 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_17_validBit[initvar] = _RAND_102[0:0];
  _RAND_105 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_17_data[initvar] = _RAND_105[3:0];
  _RAND_108 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_18_validBit[initvar] = _RAND_108[0:0];
  _RAND_111 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_18_data[initvar] = _RAND_111[3:0];
  _RAND_114 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_19_validBit[initvar] = _RAND_114[0:0];
  _RAND_117 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_19_data[initvar] = _RAND_117[3:0];
  _RAND_120 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_20_validBit[initvar] = _RAND_120[0:0];
  _RAND_123 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_20_data[initvar] = _RAND_123[3:0];
  _RAND_126 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_21_validBit[initvar] = _RAND_126[0:0];
  _RAND_129 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_21_data[initvar] = _RAND_129[3:0];
  _RAND_132 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_22_validBit[initvar] = _RAND_132[0:0];
  _RAND_135 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_22_data[initvar] = _RAND_135[3:0];
  _RAND_138 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_23_validBit[initvar] = _RAND_138[0:0];
  _RAND_141 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_23_data[initvar] = _RAND_141[3:0];
  _RAND_144 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_24_validBit[initvar] = _RAND_144[0:0];
  _RAND_147 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_24_data[initvar] = _RAND_147[3:0];
  _RAND_150 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_25_validBit[initvar] = _RAND_150[0:0];
  _RAND_153 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_25_data[initvar] = _RAND_153[3:0];
  _RAND_156 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_26_validBit[initvar] = _RAND_156[0:0];
  _RAND_159 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_26_data[initvar] = _RAND_159[3:0];
  _RAND_162 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_27_validBit[initvar] = _RAND_162[0:0];
  _RAND_165 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_27_data[initvar] = _RAND_165[3:0];
  _RAND_168 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_28_validBit[initvar] = _RAND_168[0:0];
  _RAND_171 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_28_data[initvar] = _RAND_171[3:0];
  _RAND_174 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_29_validBit[initvar] = _RAND_174[0:0];
  _RAND_177 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_29_data[initvar] = _RAND_177[3:0];
  _RAND_180 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_30_validBit[initvar] = _RAND_180[0:0];
  _RAND_183 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_30_data[initvar] = _RAND_183[3:0];
  _RAND_186 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_31_validBit[initvar] = _RAND_186[0:0];
  _RAND_189 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_31_data[initvar] = _RAND_189[3:0];
  _RAND_192 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_32_validBit[initvar] = _RAND_192[0:0];
  _RAND_195 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_32_data[initvar] = _RAND_195[3:0];
  _RAND_198 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_33_validBit[initvar] = _RAND_198[0:0];
  _RAND_201 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_33_data[initvar] = _RAND_201[3:0];
  _RAND_204 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_34_validBit[initvar] = _RAND_204[0:0];
  _RAND_207 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_34_data[initvar] = _RAND_207[3:0];
  _RAND_210 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_35_validBit[initvar] = _RAND_210[0:0];
  _RAND_213 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_35_data[initvar] = _RAND_213[3:0];
  _RAND_216 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_36_validBit[initvar] = _RAND_216[0:0];
  _RAND_219 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_36_data[initvar] = _RAND_219[3:0];
  _RAND_222 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_37_validBit[initvar] = _RAND_222[0:0];
  _RAND_225 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_37_data[initvar] = _RAND_225[3:0];
  _RAND_228 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_38_validBit[initvar] = _RAND_228[0:0];
  _RAND_231 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_38_data[initvar] = _RAND_231[3:0];
  _RAND_234 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_39_validBit[initvar] = _RAND_234[0:0];
  _RAND_237 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_39_data[initvar] = _RAND_237[3:0];
  _RAND_240 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_40_validBit[initvar] = _RAND_240[0:0];
  _RAND_243 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_40_data[initvar] = _RAND_243[3:0];
  _RAND_246 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_41_validBit[initvar] = _RAND_246[0:0];
  _RAND_249 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_41_data[initvar] = _RAND_249[3:0];
  _RAND_252 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_42_validBit[initvar] = _RAND_252[0:0];
  _RAND_255 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_42_data[initvar] = _RAND_255[3:0];
  _RAND_258 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_43_validBit[initvar] = _RAND_258[0:0];
  _RAND_261 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_43_data[initvar] = _RAND_261[3:0];
  _RAND_264 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_44_validBit[initvar] = _RAND_264[0:0];
  _RAND_267 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_44_data[initvar] = _RAND_267[3:0];
  _RAND_270 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_45_validBit[initvar] = _RAND_270[0:0];
  _RAND_273 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_45_data[initvar] = _RAND_273[3:0];
  _RAND_276 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_46_validBit[initvar] = _RAND_276[0:0];
  _RAND_279 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_46_data[initvar] = _RAND_279[3:0];
  _RAND_282 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_47_validBit[initvar] = _RAND_282[0:0];
  _RAND_285 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_47_data[initvar] = _RAND_285[3:0];
  _RAND_288 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_48_validBit[initvar] = _RAND_288[0:0];
  _RAND_291 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_48_data[initvar] = _RAND_291[3:0];
  _RAND_294 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_49_validBit[initvar] = _RAND_294[0:0];
  _RAND_297 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_49_data[initvar] = _RAND_297[3:0];
  _RAND_300 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_50_validBit[initvar] = _RAND_300[0:0];
  _RAND_303 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_50_data[initvar] = _RAND_303[3:0];
  _RAND_306 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_51_validBit[initvar] = _RAND_306[0:0];
  _RAND_309 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_51_data[initvar] = _RAND_309[3:0];
  _RAND_312 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_52_validBit[initvar] = _RAND_312[0:0];
  _RAND_315 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_52_data[initvar] = _RAND_315[3:0];
  _RAND_318 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_53_validBit[initvar] = _RAND_318[0:0];
  _RAND_321 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_53_data[initvar] = _RAND_321[3:0];
  _RAND_324 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_54_validBit[initvar] = _RAND_324[0:0];
  _RAND_327 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_54_data[initvar] = _RAND_327[3:0];
  _RAND_330 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_55_validBit[initvar] = _RAND_330[0:0];
  _RAND_333 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_55_data[initvar] = _RAND_333[3:0];
  _RAND_336 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_56_validBit[initvar] = _RAND_336[0:0];
  _RAND_339 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_56_data[initvar] = _RAND_339[3:0];
  _RAND_342 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_57_validBit[initvar] = _RAND_342[0:0];
  _RAND_345 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_57_data[initvar] = _RAND_345[3:0];
  _RAND_348 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_58_validBit[initvar] = _RAND_348[0:0];
  _RAND_351 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_58_data[initvar] = _RAND_351[3:0];
  _RAND_354 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_59_validBit[initvar] = _RAND_354[0:0];
  _RAND_357 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_59_data[initvar] = _RAND_357[3:0];
  _RAND_360 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_60_validBit[initvar] = _RAND_360[0:0];
  _RAND_363 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_60_data[initvar] = _RAND_363[3:0];
  _RAND_366 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_61_validBit[initvar] = _RAND_366[0:0];
  _RAND_369 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_61_data[initvar] = _RAND_369[3:0];
  _RAND_372 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_62_validBit[initvar] = _RAND_372[0:0];
  _RAND_375 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_62_data[initvar] = _RAND_375[3:0];
  _RAND_378 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_63_validBit[initvar] = _RAND_378[0:0];
  _RAND_381 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    inputDataBuffer_63_data[initvar] = _RAND_381[3:0];
  _RAND_384 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_0_validBit[initvar] = _RAND_384[0:0];
  _RAND_386 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_0_data[initvar] = _RAND_386[3:0];
  _RAND_388 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_1_validBit[initvar] = _RAND_388[0:0];
  _RAND_390 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_1_data[initvar] = _RAND_390[3:0];
  _RAND_392 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_2_validBit[initvar] = _RAND_392[0:0];
  _RAND_394 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_2_data[initvar] = _RAND_394[3:0];
  _RAND_396 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_3_validBit[initvar] = _RAND_396[0:0];
  _RAND_398 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_3_data[initvar] = _RAND_398[3:0];
  _RAND_400 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_4_validBit[initvar] = _RAND_400[0:0];
  _RAND_402 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_4_data[initvar] = _RAND_402[3:0];
  _RAND_404 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_5_validBit[initvar] = _RAND_404[0:0];
  _RAND_406 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_5_data[initvar] = _RAND_406[3:0];
  _RAND_408 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_6_validBit[initvar] = _RAND_408[0:0];
  _RAND_410 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_6_data[initvar] = _RAND_410[3:0];
  _RAND_412 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_7_validBit[initvar] = _RAND_412[0:0];
  _RAND_414 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_7_data[initvar] = _RAND_414[3:0];
  _RAND_416 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_8_validBit[initvar] = _RAND_416[0:0];
  _RAND_418 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_8_data[initvar] = _RAND_418[3:0];
  _RAND_420 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_9_validBit[initvar] = _RAND_420[0:0];
  _RAND_422 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_9_data[initvar] = _RAND_422[3:0];
  _RAND_424 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_10_validBit[initvar] = _RAND_424[0:0];
  _RAND_426 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_10_data[initvar] = _RAND_426[3:0];
  _RAND_428 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_11_validBit[initvar] = _RAND_428[0:0];
  _RAND_430 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_11_data[initvar] = _RAND_430[3:0];
  _RAND_432 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_12_validBit[initvar] = _RAND_432[0:0];
  _RAND_434 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_12_data[initvar] = _RAND_434[3:0];
  _RAND_436 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_13_validBit[initvar] = _RAND_436[0:0];
  _RAND_438 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_13_data[initvar] = _RAND_438[3:0];
  _RAND_440 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_14_validBit[initvar] = _RAND_440[0:0];
  _RAND_442 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_14_data[initvar] = _RAND_442[3:0];
  _RAND_444 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_15_validBit[initvar] = _RAND_444[0:0];
  _RAND_446 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_15_data[initvar] = _RAND_446[3:0];
  _RAND_448 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_16_validBit[initvar] = _RAND_448[0:0];
  _RAND_450 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_16_data[initvar] = _RAND_450[3:0];
  _RAND_452 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_17_validBit[initvar] = _RAND_452[0:0];
  _RAND_454 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_17_data[initvar] = _RAND_454[3:0];
  _RAND_456 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_18_validBit[initvar] = _RAND_456[0:0];
  _RAND_458 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_18_data[initvar] = _RAND_458[3:0];
  _RAND_460 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_19_validBit[initvar] = _RAND_460[0:0];
  _RAND_462 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_19_data[initvar] = _RAND_462[3:0];
  _RAND_464 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_20_validBit[initvar] = _RAND_464[0:0];
  _RAND_466 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_20_data[initvar] = _RAND_466[3:0];
  _RAND_468 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_21_validBit[initvar] = _RAND_468[0:0];
  _RAND_470 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_21_data[initvar] = _RAND_470[3:0];
  _RAND_472 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_22_validBit[initvar] = _RAND_472[0:0];
  _RAND_474 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_22_data[initvar] = _RAND_474[3:0];
  _RAND_476 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_23_validBit[initvar] = _RAND_476[0:0];
  _RAND_478 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_23_data[initvar] = _RAND_478[3:0];
  _RAND_480 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_24_validBit[initvar] = _RAND_480[0:0];
  _RAND_482 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_24_data[initvar] = _RAND_482[3:0];
  _RAND_484 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_25_validBit[initvar] = _RAND_484[0:0];
  _RAND_486 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_25_data[initvar] = _RAND_486[3:0];
  _RAND_488 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_26_validBit[initvar] = _RAND_488[0:0];
  _RAND_490 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_26_data[initvar] = _RAND_490[3:0];
  _RAND_492 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_27_validBit[initvar] = _RAND_492[0:0];
  _RAND_494 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_27_data[initvar] = _RAND_494[3:0];
  _RAND_496 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_28_validBit[initvar] = _RAND_496[0:0];
  _RAND_498 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_28_data[initvar] = _RAND_498[3:0];
  _RAND_500 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_29_validBit[initvar] = _RAND_500[0:0];
  _RAND_502 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_29_data[initvar] = _RAND_502[3:0];
  _RAND_504 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_30_validBit[initvar] = _RAND_504[0:0];
  _RAND_506 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_30_data[initvar] = _RAND_506[3:0];
  _RAND_508 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_31_validBit[initvar] = _RAND_508[0:0];
  _RAND_510 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_31_data[initvar] = _RAND_510[3:0];
  _RAND_512 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_32_validBit[initvar] = _RAND_512[0:0];
  _RAND_514 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_32_data[initvar] = _RAND_514[3:0];
  _RAND_516 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_33_validBit[initvar] = _RAND_516[0:0];
  _RAND_518 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_33_data[initvar] = _RAND_518[3:0];
  _RAND_520 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_34_validBit[initvar] = _RAND_520[0:0];
  _RAND_522 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_34_data[initvar] = _RAND_522[3:0];
  _RAND_524 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_35_validBit[initvar] = _RAND_524[0:0];
  _RAND_526 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_35_data[initvar] = _RAND_526[3:0];
  _RAND_528 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_36_validBit[initvar] = _RAND_528[0:0];
  _RAND_530 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_36_data[initvar] = _RAND_530[3:0];
  _RAND_532 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_37_validBit[initvar] = _RAND_532[0:0];
  _RAND_534 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_37_data[initvar] = _RAND_534[3:0];
  _RAND_536 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_38_validBit[initvar] = _RAND_536[0:0];
  _RAND_538 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_38_data[initvar] = _RAND_538[3:0];
  _RAND_540 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_39_validBit[initvar] = _RAND_540[0:0];
  _RAND_542 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_39_data[initvar] = _RAND_542[3:0];
  _RAND_544 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_40_validBit[initvar] = _RAND_544[0:0];
  _RAND_546 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_40_data[initvar] = _RAND_546[3:0];
  _RAND_548 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_41_validBit[initvar] = _RAND_548[0:0];
  _RAND_550 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_41_data[initvar] = _RAND_550[3:0];
  _RAND_552 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_42_validBit[initvar] = _RAND_552[0:0];
  _RAND_554 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_42_data[initvar] = _RAND_554[3:0];
  _RAND_556 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_43_validBit[initvar] = _RAND_556[0:0];
  _RAND_558 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_43_data[initvar] = _RAND_558[3:0];
  _RAND_560 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_44_validBit[initvar] = _RAND_560[0:0];
  _RAND_562 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_44_data[initvar] = _RAND_562[3:0];
  _RAND_564 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_45_validBit[initvar] = _RAND_564[0:0];
  _RAND_566 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_45_data[initvar] = _RAND_566[3:0];
  _RAND_568 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_46_validBit[initvar] = _RAND_568[0:0];
  _RAND_570 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_46_data[initvar] = _RAND_570[3:0];
  _RAND_572 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_47_validBit[initvar] = _RAND_572[0:0];
  _RAND_574 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_47_data[initvar] = _RAND_574[3:0];
  _RAND_576 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_48_validBit[initvar] = _RAND_576[0:0];
  _RAND_578 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_48_data[initvar] = _RAND_578[3:0];
  _RAND_580 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_49_validBit[initvar] = _RAND_580[0:0];
  _RAND_582 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_49_data[initvar] = _RAND_582[3:0];
  _RAND_584 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_50_validBit[initvar] = _RAND_584[0:0];
  _RAND_586 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_50_data[initvar] = _RAND_586[3:0];
  _RAND_588 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_51_validBit[initvar] = _RAND_588[0:0];
  _RAND_590 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_51_data[initvar] = _RAND_590[3:0];
  _RAND_592 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_52_validBit[initvar] = _RAND_592[0:0];
  _RAND_594 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_52_data[initvar] = _RAND_594[3:0];
  _RAND_596 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_53_validBit[initvar] = _RAND_596[0:0];
  _RAND_598 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_53_data[initvar] = _RAND_598[3:0];
  _RAND_600 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_54_validBit[initvar] = _RAND_600[0:0];
  _RAND_602 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_54_data[initvar] = _RAND_602[3:0];
  _RAND_604 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_55_validBit[initvar] = _RAND_604[0:0];
  _RAND_606 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_55_data[initvar] = _RAND_606[3:0];
  _RAND_608 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_56_validBit[initvar] = _RAND_608[0:0];
  _RAND_610 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_56_data[initvar] = _RAND_610[3:0];
  _RAND_612 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_57_validBit[initvar] = _RAND_612[0:0];
  _RAND_614 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_57_data[initvar] = _RAND_614[3:0];
  _RAND_616 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_58_validBit[initvar] = _RAND_616[0:0];
  _RAND_618 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_58_data[initvar] = _RAND_618[3:0];
  _RAND_620 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_59_validBit[initvar] = _RAND_620[0:0];
  _RAND_622 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_59_data[initvar] = _RAND_622[3:0];
  _RAND_624 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_60_validBit[initvar] = _RAND_624[0:0];
  _RAND_626 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_60_data[initvar] = _RAND_626[3:0];
  _RAND_628 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_61_validBit[initvar] = _RAND_628[0:0];
  _RAND_630 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_61_data[initvar] = _RAND_630[3:0];
  _RAND_632 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_62_validBit[initvar] = _RAND_632[0:0];
  _RAND_634 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_62_data[initvar] = _RAND_634[3:0];
  _RAND_636 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_63_validBit[initvar] = _RAND_636[0:0];
  _RAND_638 = {1{`RANDOM}};
  for (initvar = 0; initvar < 256; initvar = initvar+1)
    outputDataBuffer_63_data[initvar] = _RAND_638[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inputDataBuffer_0_validBit_MPORT_3_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  inputDataBuffer_0_validBit_MPORT_3_addr_pipe_0 = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  inputDataBuffer_0_data_MPORT_3_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  inputDataBuffer_0_data_MPORT_3_addr_pipe_0 = _RAND_5[7:0];
  _RAND_7 = {1{`RANDOM}};
  inputDataBuffer_1_validBit_MPORT_3_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  inputDataBuffer_1_validBit_MPORT_3_addr_pipe_0 = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  inputDataBuffer_1_data_MPORT_3_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  inputDataBuffer_1_data_MPORT_3_addr_pipe_0 = _RAND_11[7:0];
  _RAND_13 = {1{`RANDOM}};
  inputDataBuffer_2_validBit_MPORT_3_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inputDataBuffer_2_validBit_MPORT_3_addr_pipe_0 = _RAND_14[7:0];
  _RAND_16 = {1{`RANDOM}};
  inputDataBuffer_2_data_MPORT_3_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  inputDataBuffer_2_data_MPORT_3_addr_pipe_0 = _RAND_17[7:0];
  _RAND_19 = {1{`RANDOM}};
  inputDataBuffer_3_validBit_MPORT_3_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  inputDataBuffer_3_validBit_MPORT_3_addr_pipe_0 = _RAND_20[7:0];
  _RAND_22 = {1{`RANDOM}};
  inputDataBuffer_3_data_MPORT_3_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  inputDataBuffer_3_data_MPORT_3_addr_pipe_0 = _RAND_23[7:0];
  _RAND_25 = {1{`RANDOM}};
  inputDataBuffer_4_validBit_MPORT_3_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  inputDataBuffer_4_validBit_MPORT_3_addr_pipe_0 = _RAND_26[7:0];
  _RAND_28 = {1{`RANDOM}};
  inputDataBuffer_4_data_MPORT_3_en_pipe_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  inputDataBuffer_4_data_MPORT_3_addr_pipe_0 = _RAND_29[7:0];
  _RAND_31 = {1{`RANDOM}};
  inputDataBuffer_5_validBit_MPORT_3_en_pipe_0 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  inputDataBuffer_5_validBit_MPORT_3_addr_pipe_0 = _RAND_32[7:0];
  _RAND_34 = {1{`RANDOM}};
  inputDataBuffer_5_data_MPORT_3_en_pipe_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  inputDataBuffer_5_data_MPORT_3_addr_pipe_0 = _RAND_35[7:0];
  _RAND_37 = {1{`RANDOM}};
  inputDataBuffer_6_validBit_MPORT_3_en_pipe_0 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  inputDataBuffer_6_validBit_MPORT_3_addr_pipe_0 = _RAND_38[7:0];
  _RAND_40 = {1{`RANDOM}};
  inputDataBuffer_6_data_MPORT_3_en_pipe_0 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  inputDataBuffer_6_data_MPORT_3_addr_pipe_0 = _RAND_41[7:0];
  _RAND_43 = {1{`RANDOM}};
  inputDataBuffer_7_validBit_MPORT_3_en_pipe_0 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  inputDataBuffer_7_validBit_MPORT_3_addr_pipe_0 = _RAND_44[7:0];
  _RAND_46 = {1{`RANDOM}};
  inputDataBuffer_7_data_MPORT_3_en_pipe_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  inputDataBuffer_7_data_MPORT_3_addr_pipe_0 = _RAND_47[7:0];
  _RAND_49 = {1{`RANDOM}};
  inputDataBuffer_8_validBit_MPORT_3_en_pipe_0 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  inputDataBuffer_8_validBit_MPORT_3_addr_pipe_0 = _RAND_50[7:0];
  _RAND_52 = {1{`RANDOM}};
  inputDataBuffer_8_data_MPORT_3_en_pipe_0 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  inputDataBuffer_8_data_MPORT_3_addr_pipe_0 = _RAND_53[7:0];
  _RAND_55 = {1{`RANDOM}};
  inputDataBuffer_9_validBit_MPORT_3_en_pipe_0 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  inputDataBuffer_9_validBit_MPORT_3_addr_pipe_0 = _RAND_56[7:0];
  _RAND_58 = {1{`RANDOM}};
  inputDataBuffer_9_data_MPORT_3_en_pipe_0 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  inputDataBuffer_9_data_MPORT_3_addr_pipe_0 = _RAND_59[7:0];
  _RAND_61 = {1{`RANDOM}};
  inputDataBuffer_10_validBit_MPORT_3_en_pipe_0 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  inputDataBuffer_10_validBit_MPORT_3_addr_pipe_0 = _RAND_62[7:0];
  _RAND_64 = {1{`RANDOM}};
  inputDataBuffer_10_data_MPORT_3_en_pipe_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  inputDataBuffer_10_data_MPORT_3_addr_pipe_0 = _RAND_65[7:0];
  _RAND_67 = {1{`RANDOM}};
  inputDataBuffer_11_validBit_MPORT_3_en_pipe_0 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  inputDataBuffer_11_validBit_MPORT_3_addr_pipe_0 = _RAND_68[7:0];
  _RAND_70 = {1{`RANDOM}};
  inputDataBuffer_11_data_MPORT_3_en_pipe_0 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  inputDataBuffer_11_data_MPORT_3_addr_pipe_0 = _RAND_71[7:0];
  _RAND_73 = {1{`RANDOM}};
  inputDataBuffer_12_validBit_MPORT_3_en_pipe_0 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  inputDataBuffer_12_validBit_MPORT_3_addr_pipe_0 = _RAND_74[7:0];
  _RAND_76 = {1{`RANDOM}};
  inputDataBuffer_12_data_MPORT_3_en_pipe_0 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  inputDataBuffer_12_data_MPORT_3_addr_pipe_0 = _RAND_77[7:0];
  _RAND_79 = {1{`RANDOM}};
  inputDataBuffer_13_validBit_MPORT_3_en_pipe_0 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  inputDataBuffer_13_validBit_MPORT_3_addr_pipe_0 = _RAND_80[7:0];
  _RAND_82 = {1{`RANDOM}};
  inputDataBuffer_13_data_MPORT_3_en_pipe_0 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  inputDataBuffer_13_data_MPORT_3_addr_pipe_0 = _RAND_83[7:0];
  _RAND_85 = {1{`RANDOM}};
  inputDataBuffer_14_validBit_MPORT_3_en_pipe_0 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  inputDataBuffer_14_validBit_MPORT_3_addr_pipe_0 = _RAND_86[7:0];
  _RAND_88 = {1{`RANDOM}};
  inputDataBuffer_14_data_MPORT_3_en_pipe_0 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  inputDataBuffer_14_data_MPORT_3_addr_pipe_0 = _RAND_89[7:0];
  _RAND_91 = {1{`RANDOM}};
  inputDataBuffer_15_validBit_MPORT_3_en_pipe_0 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  inputDataBuffer_15_validBit_MPORT_3_addr_pipe_0 = _RAND_92[7:0];
  _RAND_94 = {1{`RANDOM}};
  inputDataBuffer_15_data_MPORT_3_en_pipe_0 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  inputDataBuffer_15_data_MPORT_3_addr_pipe_0 = _RAND_95[7:0];
  _RAND_97 = {1{`RANDOM}};
  inputDataBuffer_16_validBit_MPORT_3_en_pipe_0 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  inputDataBuffer_16_validBit_MPORT_3_addr_pipe_0 = _RAND_98[7:0];
  _RAND_100 = {1{`RANDOM}};
  inputDataBuffer_16_data_MPORT_3_en_pipe_0 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  inputDataBuffer_16_data_MPORT_3_addr_pipe_0 = _RAND_101[7:0];
  _RAND_103 = {1{`RANDOM}};
  inputDataBuffer_17_validBit_MPORT_3_en_pipe_0 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  inputDataBuffer_17_validBit_MPORT_3_addr_pipe_0 = _RAND_104[7:0];
  _RAND_106 = {1{`RANDOM}};
  inputDataBuffer_17_data_MPORT_3_en_pipe_0 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  inputDataBuffer_17_data_MPORT_3_addr_pipe_0 = _RAND_107[7:0];
  _RAND_109 = {1{`RANDOM}};
  inputDataBuffer_18_validBit_MPORT_3_en_pipe_0 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  inputDataBuffer_18_validBit_MPORT_3_addr_pipe_0 = _RAND_110[7:0];
  _RAND_112 = {1{`RANDOM}};
  inputDataBuffer_18_data_MPORT_3_en_pipe_0 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  inputDataBuffer_18_data_MPORT_3_addr_pipe_0 = _RAND_113[7:0];
  _RAND_115 = {1{`RANDOM}};
  inputDataBuffer_19_validBit_MPORT_3_en_pipe_0 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  inputDataBuffer_19_validBit_MPORT_3_addr_pipe_0 = _RAND_116[7:0];
  _RAND_118 = {1{`RANDOM}};
  inputDataBuffer_19_data_MPORT_3_en_pipe_0 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  inputDataBuffer_19_data_MPORT_3_addr_pipe_0 = _RAND_119[7:0];
  _RAND_121 = {1{`RANDOM}};
  inputDataBuffer_20_validBit_MPORT_3_en_pipe_0 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  inputDataBuffer_20_validBit_MPORT_3_addr_pipe_0 = _RAND_122[7:0];
  _RAND_124 = {1{`RANDOM}};
  inputDataBuffer_20_data_MPORT_3_en_pipe_0 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  inputDataBuffer_20_data_MPORT_3_addr_pipe_0 = _RAND_125[7:0];
  _RAND_127 = {1{`RANDOM}};
  inputDataBuffer_21_validBit_MPORT_3_en_pipe_0 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  inputDataBuffer_21_validBit_MPORT_3_addr_pipe_0 = _RAND_128[7:0];
  _RAND_130 = {1{`RANDOM}};
  inputDataBuffer_21_data_MPORT_3_en_pipe_0 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  inputDataBuffer_21_data_MPORT_3_addr_pipe_0 = _RAND_131[7:0];
  _RAND_133 = {1{`RANDOM}};
  inputDataBuffer_22_validBit_MPORT_3_en_pipe_0 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  inputDataBuffer_22_validBit_MPORT_3_addr_pipe_0 = _RAND_134[7:0];
  _RAND_136 = {1{`RANDOM}};
  inputDataBuffer_22_data_MPORT_3_en_pipe_0 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  inputDataBuffer_22_data_MPORT_3_addr_pipe_0 = _RAND_137[7:0];
  _RAND_139 = {1{`RANDOM}};
  inputDataBuffer_23_validBit_MPORT_3_en_pipe_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  inputDataBuffer_23_validBit_MPORT_3_addr_pipe_0 = _RAND_140[7:0];
  _RAND_142 = {1{`RANDOM}};
  inputDataBuffer_23_data_MPORT_3_en_pipe_0 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  inputDataBuffer_23_data_MPORT_3_addr_pipe_0 = _RAND_143[7:0];
  _RAND_145 = {1{`RANDOM}};
  inputDataBuffer_24_validBit_MPORT_3_en_pipe_0 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  inputDataBuffer_24_validBit_MPORT_3_addr_pipe_0 = _RAND_146[7:0];
  _RAND_148 = {1{`RANDOM}};
  inputDataBuffer_24_data_MPORT_3_en_pipe_0 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  inputDataBuffer_24_data_MPORT_3_addr_pipe_0 = _RAND_149[7:0];
  _RAND_151 = {1{`RANDOM}};
  inputDataBuffer_25_validBit_MPORT_3_en_pipe_0 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  inputDataBuffer_25_validBit_MPORT_3_addr_pipe_0 = _RAND_152[7:0];
  _RAND_154 = {1{`RANDOM}};
  inputDataBuffer_25_data_MPORT_3_en_pipe_0 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  inputDataBuffer_25_data_MPORT_3_addr_pipe_0 = _RAND_155[7:0];
  _RAND_157 = {1{`RANDOM}};
  inputDataBuffer_26_validBit_MPORT_3_en_pipe_0 = _RAND_157[0:0];
  _RAND_158 = {1{`RANDOM}};
  inputDataBuffer_26_validBit_MPORT_3_addr_pipe_0 = _RAND_158[7:0];
  _RAND_160 = {1{`RANDOM}};
  inputDataBuffer_26_data_MPORT_3_en_pipe_0 = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  inputDataBuffer_26_data_MPORT_3_addr_pipe_0 = _RAND_161[7:0];
  _RAND_163 = {1{`RANDOM}};
  inputDataBuffer_27_validBit_MPORT_3_en_pipe_0 = _RAND_163[0:0];
  _RAND_164 = {1{`RANDOM}};
  inputDataBuffer_27_validBit_MPORT_3_addr_pipe_0 = _RAND_164[7:0];
  _RAND_166 = {1{`RANDOM}};
  inputDataBuffer_27_data_MPORT_3_en_pipe_0 = _RAND_166[0:0];
  _RAND_167 = {1{`RANDOM}};
  inputDataBuffer_27_data_MPORT_3_addr_pipe_0 = _RAND_167[7:0];
  _RAND_169 = {1{`RANDOM}};
  inputDataBuffer_28_validBit_MPORT_3_en_pipe_0 = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  inputDataBuffer_28_validBit_MPORT_3_addr_pipe_0 = _RAND_170[7:0];
  _RAND_172 = {1{`RANDOM}};
  inputDataBuffer_28_data_MPORT_3_en_pipe_0 = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  inputDataBuffer_28_data_MPORT_3_addr_pipe_0 = _RAND_173[7:0];
  _RAND_175 = {1{`RANDOM}};
  inputDataBuffer_29_validBit_MPORT_3_en_pipe_0 = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  inputDataBuffer_29_validBit_MPORT_3_addr_pipe_0 = _RAND_176[7:0];
  _RAND_178 = {1{`RANDOM}};
  inputDataBuffer_29_data_MPORT_3_en_pipe_0 = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  inputDataBuffer_29_data_MPORT_3_addr_pipe_0 = _RAND_179[7:0];
  _RAND_181 = {1{`RANDOM}};
  inputDataBuffer_30_validBit_MPORT_3_en_pipe_0 = _RAND_181[0:0];
  _RAND_182 = {1{`RANDOM}};
  inputDataBuffer_30_validBit_MPORT_3_addr_pipe_0 = _RAND_182[7:0];
  _RAND_184 = {1{`RANDOM}};
  inputDataBuffer_30_data_MPORT_3_en_pipe_0 = _RAND_184[0:0];
  _RAND_185 = {1{`RANDOM}};
  inputDataBuffer_30_data_MPORT_3_addr_pipe_0 = _RAND_185[7:0];
  _RAND_187 = {1{`RANDOM}};
  inputDataBuffer_31_validBit_MPORT_3_en_pipe_0 = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  inputDataBuffer_31_validBit_MPORT_3_addr_pipe_0 = _RAND_188[7:0];
  _RAND_190 = {1{`RANDOM}};
  inputDataBuffer_31_data_MPORT_3_en_pipe_0 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  inputDataBuffer_31_data_MPORT_3_addr_pipe_0 = _RAND_191[7:0];
  _RAND_193 = {1{`RANDOM}};
  inputDataBuffer_32_validBit_MPORT_3_en_pipe_0 = _RAND_193[0:0];
  _RAND_194 = {1{`RANDOM}};
  inputDataBuffer_32_validBit_MPORT_3_addr_pipe_0 = _RAND_194[7:0];
  _RAND_196 = {1{`RANDOM}};
  inputDataBuffer_32_data_MPORT_3_en_pipe_0 = _RAND_196[0:0];
  _RAND_197 = {1{`RANDOM}};
  inputDataBuffer_32_data_MPORT_3_addr_pipe_0 = _RAND_197[7:0];
  _RAND_199 = {1{`RANDOM}};
  inputDataBuffer_33_validBit_MPORT_3_en_pipe_0 = _RAND_199[0:0];
  _RAND_200 = {1{`RANDOM}};
  inputDataBuffer_33_validBit_MPORT_3_addr_pipe_0 = _RAND_200[7:0];
  _RAND_202 = {1{`RANDOM}};
  inputDataBuffer_33_data_MPORT_3_en_pipe_0 = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  inputDataBuffer_33_data_MPORT_3_addr_pipe_0 = _RAND_203[7:0];
  _RAND_205 = {1{`RANDOM}};
  inputDataBuffer_34_validBit_MPORT_3_en_pipe_0 = _RAND_205[0:0];
  _RAND_206 = {1{`RANDOM}};
  inputDataBuffer_34_validBit_MPORT_3_addr_pipe_0 = _RAND_206[7:0];
  _RAND_208 = {1{`RANDOM}};
  inputDataBuffer_34_data_MPORT_3_en_pipe_0 = _RAND_208[0:0];
  _RAND_209 = {1{`RANDOM}};
  inputDataBuffer_34_data_MPORT_3_addr_pipe_0 = _RAND_209[7:0];
  _RAND_211 = {1{`RANDOM}};
  inputDataBuffer_35_validBit_MPORT_3_en_pipe_0 = _RAND_211[0:0];
  _RAND_212 = {1{`RANDOM}};
  inputDataBuffer_35_validBit_MPORT_3_addr_pipe_0 = _RAND_212[7:0];
  _RAND_214 = {1{`RANDOM}};
  inputDataBuffer_35_data_MPORT_3_en_pipe_0 = _RAND_214[0:0];
  _RAND_215 = {1{`RANDOM}};
  inputDataBuffer_35_data_MPORT_3_addr_pipe_0 = _RAND_215[7:0];
  _RAND_217 = {1{`RANDOM}};
  inputDataBuffer_36_validBit_MPORT_3_en_pipe_0 = _RAND_217[0:0];
  _RAND_218 = {1{`RANDOM}};
  inputDataBuffer_36_validBit_MPORT_3_addr_pipe_0 = _RAND_218[7:0];
  _RAND_220 = {1{`RANDOM}};
  inputDataBuffer_36_data_MPORT_3_en_pipe_0 = _RAND_220[0:0];
  _RAND_221 = {1{`RANDOM}};
  inputDataBuffer_36_data_MPORT_3_addr_pipe_0 = _RAND_221[7:0];
  _RAND_223 = {1{`RANDOM}};
  inputDataBuffer_37_validBit_MPORT_3_en_pipe_0 = _RAND_223[0:0];
  _RAND_224 = {1{`RANDOM}};
  inputDataBuffer_37_validBit_MPORT_3_addr_pipe_0 = _RAND_224[7:0];
  _RAND_226 = {1{`RANDOM}};
  inputDataBuffer_37_data_MPORT_3_en_pipe_0 = _RAND_226[0:0];
  _RAND_227 = {1{`RANDOM}};
  inputDataBuffer_37_data_MPORT_3_addr_pipe_0 = _RAND_227[7:0];
  _RAND_229 = {1{`RANDOM}};
  inputDataBuffer_38_validBit_MPORT_3_en_pipe_0 = _RAND_229[0:0];
  _RAND_230 = {1{`RANDOM}};
  inputDataBuffer_38_validBit_MPORT_3_addr_pipe_0 = _RAND_230[7:0];
  _RAND_232 = {1{`RANDOM}};
  inputDataBuffer_38_data_MPORT_3_en_pipe_0 = _RAND_232[0:0];
  _RAND_233 = {1{`RANDOM}};
  inputDataBuffer_38_data_MPORT_3_addr_pipe_0 = _RAND_233[7:0];
  _RAND_235 = {1{`RANDOM}};
  inputDataBuffer_39_validBit_MPORT_3_en_pipe_0 = _RAND_235[0:0];
  _RAND_236 = {1{`RANDOM}};
  inputDataBuffer_39_validBit_MPORT_3_addr_pipe_0 = _RAND_236[7:0];
  _RAND_238 = {1{`RANDOM}};
  inputDataBuffer_39_data_MPORT_3_en_pipe_0 = _RAND_238[0:0];
  _RAND_239 = {1{`RANDOM}};
  inputDataBuffer_39_data_MPORT_3_addr_pipe_0 = _RAND_239[7:0];
  _RAND_241 = {1{`RANDOM}};
  inputDataBuffer_40_validBit_MPORT_3_en_pipe_0 = _RAND_241[0:0];
  _RAND_242 = {1{`RANDOM}};
  inputDataBuffer_40_validBit_MPORT_3_addr_pipe_0 = _RAND_242[7:0];
  _RAND_244 = {1{`RANDOM}};
  inputDataBuffer_40_data_MPORT_3_en_pipe_0 = _RAND_244[0:0];
  _RAND_245 = {1{`RANDOM}};
  inputDataBuffer_40_data_MPORT_3_addr_pipe_0 = _RAND_245[7:0];
  _RAND_247 = {1{`RANDOM}};
  inputDataBuffer_41_validBit_MPORT_3_en_pipe_0 = _RAND_247[0:0];
  _RAND_248 = {1{`RANDOM}};
  inputDataBuffer_41_validBit_MPORT_3_addr_pipe_0 = _RAND_248[7:0];
  _RAND_250 = {1{`RANDOM}};
  inputDataBuffer_41_data_MPORT_3_en_pipe_0 = _RAND_250[0:0];
  _RAND_251 = {1{`RANDOM}};
  inputDataBuffer_41_data_MPORT_3_addr_pipe_0 = _RAND_251[7:0];
  _RAND_253 = {1{`RANDOM}};
  inputDataBuffer_42_validBit_MPORT_3_en_pipe_0 = _RAND_253[0:0];
  _RAND_254 = {1{`RANDOM}};
  inputDataBuffer_42_validBit_MPORT_3_addr_pipe_0 = _RAND_254[7:0];
  _RAND_256 = {1{`RANDOM}};
  inputDataBuffer_42_data_MPORT_3_en_pipe_0 = _RAND_256[0:0];
  _RAND_257 = {1{`RANDOM}};
  inputDataBuffer_42_data_MPORT_3_addr_pipe_0 = _RAND_257[7:0];
  _RAND_259 = {1{`RANDOM}};
  inputDataBuffer_43_validBit_MPORT_3_en_pipe_0 = _RAND_259[0:0];
  _RAND_260 = {1{`RANDOM}};
  inputDataBuffer_43_validBit_MPORT_3_addr_pipe_0 = _RAND_260[7:0];
  _RAND_262 = {1{`RANDOM}};
  inputDataBuffer_43_data_MPORT_3_en_pipe_0 = _RAND_262[0:0];
  _RAND_263 = {1{`RANDOM}};
  inputDataBuffer_43_data_MPORT_3_addr_pipe_0 = _RAND_263[7:0];
  _RAND_265 = {1{`RANDOM}};
  inputDataBuffer_44_validBit_MPORT_3_en_pipe_0 = _RAND_265[0:0];
  _RAND_266 = {1{`RANDOM}};
  inputDataBuffer_44_validBit_MPORT_3_addr_pipe_0 = _RAND_266[7:0];
  _RAND_268 = {1{`RANDOM}};
  inputDataBuffer_44_data_MPORT_3_en_pipe_0 = _RAND_268[0:0];
  _RAND_269 = {1{`RANDOM}};
  inputDataBuffer_44_data_MPORT_3_addr_pipe_0 = _RAND_269[7:0];
  _RAND_271 = {1{`RANDOM}};
  inputDataBuffer_45_validBit_MPORT_3_en_pipe_0 = _RAND_271[0:0];
  _RAND_272 = {1{`RANDOM}};
  inputDataBuffer_45_validBit_MPORT_3_addr_pipe_0 = _RAND_272[7:0];
  _RAND_274 = {1{`RANDOM}};
  inputDataBuffer_45_data_MPORT_3_en_pipe_0 = _RAND_274[0:0];
  _RAND_275 = {1{`RANDOM}};
  inputDataBuffer_45_data_MPORT_3_addr_pipe_0 = _RAND_275[7:0];
  _RAND_277 = {1{`RANDOM}};
  inputDataBuffer_46_validBit_MPORT_3_en_pipe_0 = _RAND_277[0:0];
  _RAND_278 = {1{`RANDOM}};
  inputDataBuffer_46_validBit_MPORT_3_addr_pipe_0 = _RAND_278[7:0];
  _RAND_280 = {1{`RANDOM}};
  inputDataBuffer_46_data_MPORT_3_en_pipe_0 = _RAND_280[0:0];
  _RAND_281 = {1{`RANDOM}};
  inputDataBuffer_46_data_MPORT_3_addr_pipe_0 = _RAND_281[7:0];
  _RAND_283 = {1{`RANDOM}};
  inputDataBuffer_47_validBit_MPORT_3_en_pipe_0 = _RAND_283[0:0];
  _RAND_284 = {1{`RANDOM}};
  inputDataBuffer_47_validBit_MPORT_3_addr_pipe_0 = _RAND_284[7:0];
  _RAND_286 = {1{`RANDOM}};
  inputDataBuffer_47_data_MPORT_3_en_pipe_0 = _RAND_286[0:0];
  _RAND_287 = {1{`RANDOM}};
  inputDataBuffer_47_data_MPORT_3_addr_pipe_0 = _RAND_287[7:0];
  _RAND_289 = {1{`RANDOM}};
  inputDataBuffer_48_validBit_MPORT_3_en_pipe_0 = _RAND_289[0:0];
  _RAND_290 = {1{`RANDOM}};
  inputDataBuffer_48_validBit_MPORT_3_addr_pipe_0 = _RAND_290[7:0];
  _RAND_292 = {1{`RANDOM}};
  inputDataBuffer_48_data_MPORT_3_en_pipe_0 = _RAND_292[0:0];
  _RAND_293 = {1{`RANDOM}};
  inputDataBuffer_48_data_MPORT_3_addr_pipe_0 = _RAND_293[7:0];
  _RAND_295 = {1{`RANDOM}};
  inputDataBuffer_49_validBit_MPORT_3_en_pipe_0 = _RAND_295[0:0];
  _RAND_296 = {1{`RANDOM}};
  inputDataBuffer_49_validBit_MPORT_3_addr_pipe_0 = _RAND_296[7:0];
  _RAND_298 = {1{`RANDOM}};
  inputDataBuffer_49_data_MPORT_3_en_pipe_0 = _RAND_298[0:0];
  _RAND_299 = {1{`RANDOM}};
  inputDataBuffer_49_data_MPORT_3_addr_pipe_0 = _RAND_299[7:0];
  _RAND_301 = {1{`RANDOM}};
  inputDataBuffer_50_validBit_MPORT_3_en_pipe_0 = _RAND_301[0:0];
  _RAND_302 = {1{`RANDOM}};
  inputDataBuffer_50_validBit_MPORT_3_addr_pipe_0 = _RAND_302[7:0];
  _RAND_304 = {1{`RANDOM}};
  inputDataBuffer_50_data_MPORT_3_en_pipe_0 = _RAND_304[0:0];
  _RAND_305 = {1{`RANDOM}};
  inputDataBuffer_50_data_MPORT_3_addr_pipe_0 = _RAND_305[7:0];
  _RAND_307 = {1{`RANDOM}};
  inputDataBuffer_51_validBit_MPORT_3_en_pipe_0 = _RAND_307[0:0];
  _RAND_308 = {1{`RANDOM}};
  inputDataBuffer_51_validBit_MPORT_3_addr_pipe_0 = _RAND_308[7:0];
  _RAND_310 = {1{`RANDOM}};
  inputDataBuffer_51_data_MPORT_3_en_pipe_0 = _RAND_310[0:0];
  _RAND_311 = {1{`RANDOM}};
  inputDataBuffer_51_data_MPORT_3_addr_pipe_0 = _RAND_311[7:0];
  _RAND_313 = {1{`RANDOM}};
  inputDataBuffer_52_validBit_MPORT_3_en_pipe_0 = _RAND_313[0:0];
  _RAND_314 = {1{`RANDOM}};
  inputDataBuffer_52_validBit_MPORT_3_addr_pipe_0 = _RAND_314[7:0];
  _RAND_316 = {1{`RANDOM}};
  inputDataBuffer_52_data_MPORT_3_en_pipe_0 = _RAND_316[0:0];
  _RAND_317 = {1{`RANDOM}};
  inputDataBuffer_52_data_MPORT_3_addr_pipe_0 = _RAND_317[7:0];
  _RAND_319 = {1{`RANDOM}};
  inputDataBuffer_53_validBit_MPORT_3_en_pipe_0 = _RAND_319[0:0];
  _RAND_320 = {1{`RANDOM}};
  inputDataBuffer_53_validBit_MPORT_3_addr_pipe_0 = _RAND_320[7:0];
  _RAND_322 = {1{`RANDOM}};
  inputDataBuffer_53_data_MPORT_3_en_pipe_0 = _RAND_322[0:0];
  _RAND_323 = {1{`RANDOM}};
  inputDataBuffer_53_data_MPORT_3_addr_pipe_0 = _RAND_323[7:0];
  _RAND_325 = {1{`RANDOM}};
  inputDataBuffer_54_validBit_MPORT_3_en_pipe_0 = _RAND_325[0:0];
  _RAND_326 = {1{`RANDOM}};
  inputDataBuffer_54_validBit_MPORT_3_addr_pipe_0 = _RAND_326[7:0];
  _RAND_328 = {1{`RANDOM}};
  inputDataBuffer_54_data_MPORT_3_en_pipe_0 = _RAND_328[0:0];
  _RAND_329 = {1{`RANDOM}};
  inputDataBuffer_54_data_MPORT_3_addr_pipe_0 = _RAND_329[7:0];
  _RAND_331 = {1{`RANDOM}};
  inputDataBuffer_55_validBit_MPORT_3_en_pipe_0 = _RAND_331[0:0];
  _RAND_332 = {1{`RANDOM}};
  inputDataBuffer_55_validBit_MPORT_3_addr_pipe_0 = _RAND_332[7:0];
  _RAND_334 = {1{`RANDOM}};
  inputDataBuffer_55_data_MPORT_3_en_pipe_0 = _RAND_334[0:0];
  _RAND_335 = {1{`RANDOM}};
  inputDataBuffer_55_data_MPORT_3_addr_pipe_0 = _RAND_335[7:0];
  _RAND_337 = {1{`RANDOM}};
  inputDataBuffer_56_validBit_MPORT_3_en_pipe_0 = _RAND_337[0:0];
  _RAND_338 = {1{`RANDOM}};
  inputDataBuffer_56_validBit_MPORT_3_addr_pipe_0 = _RAND_338[7:0];
  _RAND_340 = {1{`RANDOM}};
  inputDataBuffer_56_data_MPORT_3_en_pipe_0 = _RAND_340[0:0];
  _RAND_341 = {1{`RANDOM}};
  inputDataBuffer_56_data_MPORT_3_addr_pipe_0 = _RAND_341[7:0];
  _RAND_343 = {1{`RANDOM}};
  inputDataBuffer_57_validBit_MPORT_3_en_pipe_0 = _RAND_343[0:0];
  _RAND_344 = {1{`RANDOM}};
  inputDataBuffer_57_validBit_MPORT_3_addr_pipe_0 = _RAND_344[7:0];
  _RAND_346 = {1{`RANDOM}};
  inputDataBuffer_57_data_MPORT_3_en_pipe_0 = _RAND_346[0:0];
  _RAND_347 = {1{`RANDOM}};
  inputDataBuffer_57_data_MPORT_3_addr_pipe_0 = _RAND_347[7:0];
  _RAND_349 = {1{`RANDOM}};
  inputDataBuffer_58_validBit_MPORT_3_en_pipe_0 = _RAND_349[0:0];
  _RAND_350 = {1{`RANDOM}};
  inputDataBuffer_58_validBit_MPORT_3_addr_pipe_0 = _RAND_350[7:0];
  _RAND_352 = {1{`RANDOM}};
  inputDataBuffer_58_data_MPORT_3_en_pipe_0 = _RAND_352[0:0];
  _RAND_353 = {1{`RANDOM}};
  inputDataBuffer_58_data_MPORT_3_addr_pipe_0 = _RAND_353[7:0];
  _RAND_355 = {1{`RANDOM}};
  inputDataBuffer_59_validBit_MPORT_3_en_pipe_0 = _RAND_355[0:0];
  _RAND_356 = {1{`RANDOM}};
  inputDataBuffer_59_validBit_MPORT_3_addr_pipe_0 = _RAND_356[7:0];
  _RAND_358 = {1{`RANDOM}};
  inputDataBuffer_59_data_MPORT_3_en_pipe_0 = _RAND_358[0:0];
  _RAND_359 = {1{`RANDOM}};
  inputDataBuffer_59_data_MPORT_3_addr_pipe_0 = _RAND_359[7:0];
  _RAND_361 = {1{`RANDOM}};
  inputDataBuffer_60_validBit_MPORT_3_en_pipe_0 = _RAND_361[0:0];
  _RAND_362 = {1{`RANDOM}};
  inputDataBuffer_60_validBit_MPORT_3_addr_pipe_0 = _RAND_362[7:0];
  _RAND_364 = {1{`RANDOM}};
  inputDataBuffer_60_data_MPORT_3_en_pipe_0 = _RAND_364[0:0];
  _RAND_365 = {1{`RANDOM}};
  inputDataBuffer_60_data_MPORT_3_addr_pipe_0 = _RAND_365[7:0];
  _RAND_367 = {1{`RANDOM}};
  inputDataBuffer_61_validBit_MPORT_3_en_pipe_0 = _RAND_367[0:0];
  _RAND_368 = {1{`RANDOM}};
  inputDataBuffer_61_validBit_MPORT_3_addr_pipe_0 = _RAND_368[7:0];
  _RAND_370 = {1{`RANDOM}};
  inputDataBuffer_61_data_MPORT_3_en_pipe_0 = _RAND_370[0:0];
  _RAND_371 = {1{`RANDOM}};
  inputDataBuffer_61_data_MPORT_3_addr_pipe_0 = _RAND_371[7:0];
  _RAND_373 = {1{`RANDOM}};
  inputDataBuffer_62_validBit_MPORT_3_en_pipe_0 = _RAND_373[0:0];
  _RAND_374 = {1{`RANDOM}};
  inputDataBuffer_62_validBit_MPORT_3_addr_pipe_0 = _RAND_374[7:0];
  _RAND_376 = {1{`RANDOM}};
  inputDataBuffer_62_data_MPORT_3_en_pipe_0 = _RAND_376[0:0];
  _RAND_377 = {1{`RANDOM}};
  inputDataBuffer_62_data_MPORT_3_addr_pipe_0 = _RAND_377[7:0];
  _RAND_379 = {1{`RANDOM}};
  inputDataBuffer_63_validBit_MPORT_3_en_pipe_0 = _RAND_379[0:0];
  _RAND_380 = {1{`RANDOM}};
  inputDataBuffer_63_validBit_MPORT_3_addr_pipe_0 = _RAND_380[7:0];
  _RAND_382 = {1{`RANDOM}};
  inputDataBuffer_63_data_MPORT_3_en_pipe_0 = _RAND_382[0:0];
  _RAND_383 = {1{`RANDOM}};
  inputDataBuffer_63_data_MPORT_3_addr_pipe_0 = _RAND_383[7:0];
  _RAND_385 = {1{`RANDOM}};
  outputDataBuffer_0_validBit_MPORT_2_addr_pipe_0 = _RAND_385[7:0];
  _RAND_387 = {1{`RANDOM}};
  outputDataBuffer_0_data_MPORT_2_addr_pipe_0 = _RAND_387[7:0];
  _RAND_389 = {1{`RANDOM}};
  outputDataBuffer_1_validBit_MPORT_2_addr_pipe_0 = _RAND_389[7:0];
  _RAND_391 = {1{`RANDOM}};
  outputDataBuffer_1_data_MPORT_2_addr_pipe_0 = _RAND_391[7:0];
  _RAND_393 = {1{`RANDOM}};
  outputDataBuffer_2_validBit_MPORT_2_addr_pipe_0 = _RAND_393[7:0];
  _RAND_395 = {1{`RANDOM}};
  outputDataBuffer_2_data_MPORT_2_addr_pipe_0 = _RAND_395[7:0];
  _RAND_397 = {1{`RANDOM}};
  outputDataBuffer_3_validBit_MPORT_2_addr_pipe_0 = _RAND_397[7:0];
  _RAND_399 = {1{`RANDOM}};
  outputDataBuffer_3_data_MPORT_2_addr_pipe_0 = _RAND_399[7:0];
  _RAND_401 = {1{`RANDOM}};
  outputDataBuffer_4_validBit_MPORT_2_addr_pipe_0 = _RAND_401[7:0];
  _RAND_403 = {1{`RANDOM}};
  outputDataBuffer_4_data_MPORT_2_addr_pipe_0 = _RAND_403[7:0];
  _RAND_405 = {1{`RANDOM}};
  outputDataBuffer_5_validBit_MPORT_2_addr_pipe_0 = _RAND_405[7:0];
  _RAND_407 = {1{`RANDOM}};
  outputDataBuffer_5_data_MPORT_2_addr_pipe_0 = _RAND_407[7:0];
  _RAND_409 = {1{`RANDOM}};
  outputDataBuffer_6_validBit_MPORT_2_addr_pipe_0 = _RAND_409[7:0];
  _RAND_411 = {1{`RANDOM}};
  outputDataBuffer_6_data_MPORT_2_addr_pipe_0 = _RAND_411[7:0];
  _RAND_413 = {1{`RANDOM}};
  outputDataBuffer_7_validBit_MPORT_2_addr_pipe_0 = _RAND_413[7:0];
  _RAND_415 = {1{`RANDOM}};
  outputDataBuffer_7_data_MPORT_2_addr_pipe_0 = _RAND_415[7:0];
  _RAND_417 = {1{`RANDOM}};
  outputDataBuffer_8_validBit_MPORT_2_addr_pipe_0 = _RAND_417[7:0];
  _RAND_419 = {1{`RANDOM}};
  outputDataBuffer_8_data_MPORT_2_addr_pipe_0 = _RAND_419[7:0];
  _RAND_421 = {1{`RANDOM}};
  outputDataBuffer_9_validBit_MPORT_2_addr_pipe_0 = _RAND_421[7:0];
  _RAND_423 = {1{`RANDOM}};
  outputDataBuffer_9_data_MPORT_2_addr_pipe_0 = _RAND_423[7:0];
  _RAND_425 = {1{`RANDOM}};
  outputDataBuffer_10_validBit_MPORT_2_addr_pipe_0 = _RAND_425[7:0];
  _RAND_427 = {1{`RANDOM}};
  outputDataBuffer_10_data_MPORT_2_addr_pipe_0 = _RAND_427[7:0];
  _RAND_429 = {1{`RANDOM}};
  outputDataBuffer_11_validBit_MPORT_2_addr_pipe_0 = _RAND_429[7:0];
  _RAND_431 = {1{`RANDOM}};
  outputDataBuffer_11_data_MPORT_2_addr_pipe_0 = _RAND_431[7:0];
  _RAND_433 = {1{`RANDOM}};
  outputDataBuffer_12_validBit_MPORT_2_addr_pipe_0 = _RAND_433[7:0];
  _RAND_435 = {1{`RANDOM}};
  outputDataBuffer_12_data_MPORT_2_addr_pipe_0 = _RAND_435[7:0];
  _RAND_437 = {1{`RANDOM}};
  outputDataBuffer_13_validBit_MPORT_2_addr_pipe_0 = _RAND_437[7:0];
  _RAND_439 = {1{`RANDOM}};
  outputDataBuffer_13_data_MPORT_2_addr_pipe_0 = _RAND_439[7:0];
  _RAND_441 = {1{`RANDOM}};
  outputDataBuffer_14_validBit_MPORT_2_addr_pipe_0 = _RAND_441[7:0];
  _RAND_443 = {1{`RANDOM}};
  outputDataBuffer_14_data_MPORT_2_addr_pipe_0 = _RAND_443[7:0];
  _RAND_445 = {1{`RANDOM}};
  outputDataBuffer_15_validBit_MPORT_2_addr_pipe_0 = _RAND_445[7:0];
  _RAND_447 = {1{`RANDOM}};
  outputDataBuffer_15_data_MPORT_2_addr_pipe_0 = _RAND_447[7:0];
  _RAND_449 = {1{`RANDOM}};
  outputDataBuffer_16_validBit_MPORT_2_addr_pipe_0 = _RAND_449[7:0];
  _RAND_451 = {1{`RANDOM}};
  outputDataBuffer_16_data_MPORT_2_addr_pipe_0 = _RAND_451[7:0];
  _RAND_453 = {1{`RANDOM}};
  outputDataBuffer_17_validBit_MPORT_2_addr_pipe_0 = _RAND_453[7:0];
  _RAND_455 = {1{`RANDOM}};
  outputDataBuffer_17_data_MPORT_2_addr_pipe_0 = _RAND_455[7:0];
  _RAND_457 = {1{`RANDOM}};
  outputDataBuffer_18_validBit_MPORT_2_addr_pipe_0 = _RAND_457[7:0];
  _RAND_459 = {1{`RANDOM}};
  outputDataBuffer_18_data_MPORT_2_addr_pipe_0 = _RAND_459[7:0];
  _RAND_461 = {1{`RANDOM}};
  outputDataBuffer_19_validBit_MPORT_2_addr_pipe_0 = _RAND_461[7:0];
  _RAND_463 = {1{`RANDOM}};
  outputDataBuffer_19_data_MPORT_2_addr_pipe_0 = _RAND_463[7:0];
  _RAND_465 = {1{`RANDOM}};
  outputDataBuffer_20_validBit_MPORT_2_addr_pipe_0 = _RAND_465[7:0];
  _RAND_467 = {1{`RANDOM}};
  outputDataBuffer_20_data_MPORT_2_addr_pipe_0 = _RAND_467[7:0];
  _RAND_469 = {1{`RANDOM}};
  outputDataBuffer_21_validBit_MPORT_2_addr_pipe_0 = _RAND_469[7:0];
  _RAND_471 = {1{`RANDOM}};
  outputDataBuffer_21_data_MPORT_2_addr_pipe_0 = _RAND_471[7:0];
  _RAND_473 = {1{`RANDOM}};
  outputDataBuffer_22_validBit_MPORT_2_addr_pipe_0 = _RAND_473[7:0];
  _RAND_475 = {1{`RANDOM}};
  outputDataBuffer_22_data_MPORT_2_addr_pipe_0 = _RAND_475[7:0];
  _RAND_477 = {1{`RANDOM}};
  outputDataBuffer_23_validBit_MPORT_2_addr_pipe_0 = _RAND_477[7:0];
  _RAND_479 = {1{`RANDOM}};
  outputDataBuffer_23_data_MPORT_2_addr_pipe_0 = _RAND_479[7:0];
  _RAND_481 = {1{`RANDOM}};
  outputDataBuffer_24_validBit_MPORT_2_addr_pipe_0 = _RAND_481[7:0];
  _RAND_483 = {1{`RANDOM}};
  outputDataBuffer_24_data_MPORT_2_addr_pipe_0 = _RAND_483[7:0];
  _RAND_485 = {1{`RANDOM}};
  outputDataBuffer_25_validBit_MPORT_2_addr_pipe_0 = _RAND_485[7:0];
  _RAND_487 = {1{`RANDOM}};
  outputDataBuffer_25_data_MPORT_2_addr_pipe_0 = _RAND_487[7:0];
  _RAND_489 = {1{`RANDOM}};
  outputDataBuffer_26_validBit_MPORT_2_addr_pipe_0 = _RAND_489[7:0];
  _RAND_491 = {1{`RANDOM}};
  outputDataBuffer_26_data_MPORT_2_addr_pipe_0 = _RAND_491[7:0];
  _RAND_493 = {1{`RANDOM}};
  outputDataBuffer_27_validBit_MPORT_2_addr_pipe_0 = _RAND_493[7:0];
  _RAND_495 = {1{`RANDOM}};
  outputDataBuffer_27_data_MPORT_2_addr_pipe_0 = _RAND_495[7:0];
  _RAND_497 = {1{`RANDOM}};
  outputDataBuffer_28_validBit_MPORT_2_addr_pipe_0 = _RAND_497[7:0];
  _RAND_499 = {1{`RANDOM}};
  outputDataBuffer_28_data_MPORT_2_addr_pipe_0 = _RAND_499[7:0];
  _RAND_501 = {1{`RANDOM}};
  outputDataBuffer_29_validBit_MPORT_2_addr_pipe_0 = _RAND_501[7:0];
  _RAND_503 = {1{`RANDOM}};
  outputDataBuffer_29_data_MPORT_2_addr_pipe_0 = _RAND_503[7:0];
  _RAND_505 = {1{`RANDOM}};
  outputDataBuffer_30_validBit_MPORT_2_addr_pipe_0 = _RAND_505[7:0];
  _RAND_507 = {1{`RANDOM}};
  outputDataBuffer_30_data_MPORT_2_addr_pipe_0 = _RAND_507[7:0];
  _RAND_509 = {1{`RANDOM}};
  outputDataBuffer_31_validBit_MPORT_2_addr_pipe_0 = _RAND_509[7:0];
  _RAND_511 = {1{`RANDOM}};
  outputDataBuffer_31_data_MPORT_2_addr_pipe_0 = _RAND_511[7:0];
  _RAND_513 = {1{`RANDOM}};
  outputDataBuffer_32_validBit_MPORT_2_addr_pipe_0 = _RAND_513[7:0];
  _RAND_515 = {1{`RANDOM}};
  outputDataBuffer_32_data_MPORT_2_addr_pipe_0 = _RAND_515[7:0];
  _RAND_517 = {1{`RANDOM}};
  outputDataBuffer_33_validBit_MPORT_2_addr_pipe_0 = _RAND_517[7:0];
  _RAND_519 = {1{`RANDOM}};
  outputDataBuffer_33_data_MPORT_2_addr_pipe_0 = _RAND_519[7:0];
  _RAND_521 = {1{`RANDOM}};
  outputDataBuffer_34_validBit_MPORT_2_addr_pipe_0 = _RAND_521[7:0];
  _RAND_523 = {1{`RANDOM}};
  outputDataBuffer_34_data_MPORT_2_addr_pipe_0 = _RAND_523[7:0];
  _RAND_525 = {1{`RANDOM}};
  outputDataBuffer_35_validBit_MPORT_2_addr_pipe_0 = _RAND_525[7:0];
  _RAND_527 = {1{`RANDOM}};
  outputDataBuffer_35_data_MPORT_2_addr_pipe_0 = _RAND_527[7:0];
  _RAND_529 = {1{`RANDOM}};
  outputDataBuffer_36_validBit_MPORT_2_addr_pipe_0 = _RAND_529[7:0];
  _RAND_531 = {1{`RANDOM}};
  outputDataBuffer_36_data_MPORT_2_addr_pipe_0 = _RAND_531[7:0];
  _RAND_533 = {1{`RANDOM}};
  outputDataBuffer_37_validBit_MPORT_2_addr_pipe_0 = _RAND_533[7:0];
  _RAND_535 = {1{`RANDOM}};
  outputDataBuffer_37_data_MPORT_2_addr_pipe_0 = _RAND_535[7:0];
  _RAND_537 = {1{`RANDOM}};
  outputDataBuffer_38_validBit_MPORT_2_addr_pipe_0 = _RAND_537[7:0];
  _RAND_539 = {1{`RANDOM}};
  outputDataBuffer_38_data_MPORT_2_addr_pipe_0 = _RAND_539[7:0];
  _RAND_541 = {1{`RANDOM}};
  outputDataBuffer_39_validBit_MPORT_2_addr_pipe_0 = _RAND_541[7:0];
  _RAND_543 = {1{`RANDOM}};
  outputDataBuffer_39_data_MPORT_2_addr_pipe_0 = _RAND_543[7:0];
  _RAND_545 = {1{`RANDOM}};
  outputDataBuffer_40_validBit_MPORT_2_addr_pipe_0 = _RAND_545[7:0];
  _RAND_547 = {1{`RANDOM}};
  outputDataBuffer_40_data_MPORT_2_addr_pipe_0 = _RAND_547[7:0];
  _RAND_549 = {1{`RANDOM}};
  outputDataBuffer_41_validBit_MPORT_2_addr_pipe_0 = _RAND_549[7:0];
  _RAND_551 = {1{`RANDOM}};
  outputDataBuffer_41_data_MPORT_2_addr_pipe_0 = _RAND_551[7:0];
  _RAND_553 = {1{`RANDOM}};
  outputDataBuffer_42_validBit_MPORT_2_addr_pipe_0 = _RAND_553[7:0];
  _RAND_555 = {1{`RANDOM}};
  outputDataBuffer_42_data_MPORT_2_addr_pipe_0 = _RAND_555[7:0];
  _RAND_557 = {1{`RANDOM}};
  outputDataBuffer_43_validBit_MPORT_2_addr_pipe_0 = _RAND_557[7:0];
  _RAND_559 = {1{`RANDOM}};
  outputDataBuffer_43_data_MPORT_2_addr_pipe_0 = _RAND_559[7:0];
  _RAND_561 = {1{`RANDOM}};
  outputDataBuffer_44_validBit_MPORT_2_addr_pipe_0 = _RAND_561[7:0];
  _RAND_563 = {1{`RANDOM}};
  outputDataBuffer_44_data_MPORT_2_addr_pipe_0 = _RAND_563[7:0];
  _RAND_565 = {1{`RANDOM}};
  outputDataBuffer_45_validBit_MPORT_2_addr_pipe_0 = _RAND_565[7:0];
  _RAND_567 = {1{`RANDOM}};
  outputDataBuffer_45_data_MPORT_2_addr_pipe_0 = _RAND_567[7:0];
  _RAND_569 = {1{`RANDOM}};
  outputDataBuffer_46_validBit_MPORT_2_addr_pipe_0 = _RAND_569[7:0];
  _RAND_571 = {1{`RANDOM}};
  outputDataBuffer_46_data_MPORT_2_addr_pipe_0 = _RAND_571[7:0];
  _RAND_573 = {1{`RANDOM}};
  outputDataBuffer_47_validBit_MPORT_2_addr_pipe_0 = _RAND_573[7:0];
  _RAND_575 = {1{`RANDOM}};
  outputDataBuffer_47_data_MPORT_2_addr_pipe_0 = _RAND_575[7:0];
  _RAND_577 = {1{`RANDOM}};
  outputDataBuffer_48_validBit_MPORT_2_addr_pipe_0 = _RAND_577[7:0];
  _RAND_579 = {1{`RANDOM}};
  outputDataBuffer_48_data_MPORT_2_addr_pipe_0 = _RAND_579[7:0];
  _RAND_581 = {1{`RANDOM}};
  outputDataBuffer_49_validBit_MPORT_2_addr_pipe_0 = _RAND_581[7:0];
  _RAND_583 = {1{`RANDOM}};
  outputDataBuffer_49_data_MPORT_2_addr_pipe_0 = _RAND_583[7:0];
  _RAND_585 = {1{`RANDOM}};
  outputDataBuffer_50_validBit_MPORT_2_addr_pipe_0 = _RAND_585[7:0];
  _RAND_587 = {1{`RANDOM}};
  outputDataBuffer_50_data_MPORT_2_addr_pipe_0 = _RAND_587[7:0];
  _RAND_589 = {1{`RANDOM}};
  outputDataBuffer_51_validBit_MPORT_2_addr_pipe_0 = _RAND_589[7:0];
  _RAND_591 = {1{`RANDOM}};
  outputDataBuffer_51_data_MPORT_2_addr_pipe_0 = _RAND_591[7:0];
  _RAND_593 = {1{`RANDOM}};
  outputDataBuffer_52_validBit_MPORT_2_addr_pipe_0 = _RAND_593[7:0];
  _RAND_595 = {1{`RANDOM}};
  outputDataBuffer_52_data_MPORT_2_addr_pipe_0 = _RAND_595[7:0];
  _RAND_597 = {1{`RANDOM}};
  outputDataBuffer_53_validBit_MPORT_2_addr_pipe_0 = _RAND_597[7:0];
  _RAND_599 = {1{`RANDOM}};
  outputDataBuffer_53_data_MPORT_2_addr_pipe_0 = _RAND_599[7:0];
  _RAND_601 = {1{`RANDOM}};
  outputDataBuffer_54_validBit_MPORT_2_addr_pipe_0 = _RAND_601[7:0];
  _RAND_603 = {1{`RANDOM}};
  outputDataBuffer_54_data_MPORT_2_addr_pipe_0 = _RAND_603[7:0];
  _RAND_605 = {1{`RANDOM}};
  outputDataBuffer_55_validBit_MPORT_2_addr_pipe_0 = _RAND_605[7:0];
  _RAND_607 = {1{`RANDOM}};
  outputDataBuffer_55_data_MPORT_2_addr_pipe_0 = _RAND_607[7:0];
  _RAND_609 = {1{`RANDOM}};
  outputDataBuffer_56_validBit_MPORT_2_addr_pipe_0 = _RAND_609[7:0];
  _RAND_611 = {1{`RANDOM}};
  outputDataBuffer_56_data_MPORT_2_addr_pipe_0 = _RAND_611[7:0];
  _RAND_613 = {1{`RANDOM}};
  outputDataBuffer_57_validBit_MPORT_2_addr_pipe_0 = _RAND_613[7:0];
  _RAND_615 = {1{`RANDOM}};
  outputDataBuffer_57_data_MPORT_2_addr_pipe_0 = _RAND_615[7:0];
  _RAND_617 = {1{`RANDOM}};
  outputDataBuffer_58_validBit_MPORT_2_addr_pipe_0 = _RAND_617[7:0];
  _RAND_619 = {1{`RANDOM}};
  outputDataBuffer_58_data_MPORT_2_addr_pipe_0 = _RAND_619[7:0];
  _RAND_621 = {1{`RANDOM}};
  outputDataBuffer_59_validBit_MPORT_2_addr_pipe_0 = _RAND_621[7:0];
  _RAND_623 = {1{`RANDOM}};
  outputDataBuffer_59_data_MPORT_2_addr_pipe_0 = _RAND_623[7:0];
  _RAND_625 = {1{`RANDOM}};
  outputDataBuffer_60_validBit_MPORT_2_addr_pipe_0 = _RAND_625[7:0];
  _RAND_627 = {1{`RANDOM}};
  outputDataBuffer_60_data_MPORT_2_addr_pipe_0 = _RAND_627[7:0];
  _RAND_629 = {1{`RANDOM}};
  outputDataBuffer_61_validBit_MPORT_2_addr_pipe_0 = _RAND_629[7:0];
  _RAND_631 = {1{`RANDOM}};
  outputDataBuffer_61_data_MPORT_2_addr_pipe_0 = _RAND_631[7:0];
  _RAND_633 = {1{`RANDOM}};
  outputDataBuffer_62_validBit_MPORT_2_addr_pipe_0 = _RAND_633[7:0];
  _RAND_635 = {1{`RANDOM}};
  outputDataBuffer_62_data_MPORT_2_addr_pipe_0 = _RAND_635[7:0];
  _RAND_637 = {1{`RANDOM}};
  outputDataBuffer_63_validBit_MPORT_2_addr_pipe_0 = _RAND_637[7:0];
  _RAND_639 = {1{`RANDOM}};
  outputDataBuffer_63_data_MPORT_2_addr_pipe_0 = _RAND_639[7:0];
  _RAND_640 = {1{`RANDOM}};
  wr_Addr_inBuf = _RAND_640[7:0];
  _RAND_641 = {1{`RANDOM}};
  rd_Addr_inBuf = _RAND_641[7:0];
  _RAND_642 = {1{`RANDOM}};
  rd_D_inBuf_0_validBit = _RAND_642[0:0];
  _RAND_643 = {1{`RANDOM}};
  rd_D_inBuf_0_data = _RAND_643[3:0];
  _RAND_644 = {1{`RANDOM}};
  rd_D_inBuf_1_validBit = _RAND_644[0:0];
  _RAND_645 = {1{`RANDOM}};
  rd_D_inBuf_1_data = _RAND_645[3:0];
  _RAND_646 = {1{`RANDOM}};
  rd_D_inBuf_2_validBit = _RAND_646[0:0];
  _RAND_647 = {1{`RANDOM}};
  rd_D_inBuf_2_data = _RAND_647[3:0];
  _RAND_648 = {1{`RANDOM}};
  rd_D_inBuf_3_validBit = _RAND_648[0:0];
  _RAND_649 = {1{`RANDOM}};
  rd_D_inBuf_3_data = _RAND_649[3:0];
  _RAND_650 = {1{`RANDOM}};
  rd_D_inBuf_4_validBit = _RAND_650[0:0];
  _RAND_651 = {1{`RANDOM}};
  rd_D_inBuf_4_data = _RAND_651[3:0];
  _RAND_652 = {1{`RANDOM}};
  rd_D_inBuf_5_validBit = _RAND_652[0:0];
  _RAND_653 = {1{`RANDOM}};
  rd_D_inBuf_5_data = _RAND_653[3:0];
  _RAND_654 = {1{`RANDOM}};
  rd_D_inBuf_6_validBit = _RAND_654[0:0];
  _RAND_655 = {1{`RANDOM}};
  rd_D_inBuf_6_data = _RAND_655[3:0];
  _RAND_656 = {1{`RANDOM}};
  rd_D_inBuf_7_validBit = _RAND_656[0:0];
  _RAND_657 = {1{`RANDOM}};
  rd_D_inBuf_7_data = _RAND_657[3:0];
  _RAND_658 = {1{`RANDOM}};
  rd_D_inBuf_8_validBit = _RAND_658[0:0];
  _RAND_659 = {1{`RANDOM}};
  rd_D_inBuf_8_data = _RAND_659[3:0];
  _RAND_660 = {1{`RANDOM}};
  rd_D_inBuf_9_validBit = _RAND_660[0:0];
  _RAND_661 = {1{`RANDOM}};
  rd_D_inBuf_9_data = _RAND_661[3:0];
  _RAND_662 = {1{`RANDOM}};
  rd_D_inBuf_10_validBit = _RAND_662[0:0];
  _RAND_663 = {1{`RANDOM}};
  rd_D_inBuf_10_data = _RAND_663[3:0];
  _RAND_664 = {1{`RANDOM}};
  rd_D_inBuf_11_validBit = _RAND_664[0:0];
  _RAND_665 = {1{`RANDOM}};
  rd_D_inBuf_11_data = _RAND_665[3:0];
  _RAND_666 = {1{`RANDOM}};
  rd_D_inBuf_12_validBit = _RAND_666[0:0];
  _RAND_667 = {1{`RANDOM}};
  rd_D_inBuf_12_data = _RAND_667[3:0];
  _RAND_668 = {1{`RANDOM}};
  rd_D_inBuf_13_validBit = _RAND_668[0:0];
  _RAND_669 = {1{`RANDOM}};
  rd_D_inBuf_13_data = _RAND_669[3:0];
  _RAND_670 = {1{`RANDOM}};
  rd_D_inBuf_14_validBit = _RAND_670[0:0];
  _RAND_671 = {1{`RANDOM}};
  rd_D_inBuf_14_data = _RAND_671[3:0];
  _RAND_672 = {1{`RANDOM}};
  rd_D_inBuf_15_validBit = _RAND_672[0:0];
  _RAND_673 = {1{`RANDOM}};
  rd_D_inBuf_15_data = _RAND_673[3:0];
  _RAND_674 = {1{`RANDOM}};
  rd_D_inBuf_16_validBit = _RAND_674[0:0];
  _RAND_675 = {1{`RANDOM}};
  rd_D_inBuf_16_data = _RAND_675[3:0];
  _RAND_676 = {1{`RANDOM}};
  rd_D_inBuf_17_validBit = _RAND_676[0:0];
  _RAND_677 = {1{`RANDOM}};
  rd_D_inBuf_17_data = _RAND_677[3:0];
  _RAND_678 = {1{`RANDOM}};
  rd_D_inBuf_18_validBit = _RAND_678[0:0];
  _RAND_679 = {1{`RANDOM}};
  rd_D_inBuf_18_data = _RAND_679[3:0];
  _RAND_680 = {1{`RANDOM}};
  rd_D_inBuf_19_validBit = _RAND_680[0:0];
  _RAND_681 = {1{`RANDOM}};
  rd_D_inBuf_19_data = _RAND_681[3:0];
  _RAND_682 = {1{`RANDOM}};
  rd_D_inBuf_20_validBit = _RAND_682[0:0];
  _RAND_683 = {1{`RANDOM}};
  rd_D_inBuf_20_data = _RAND_683[3:0];
  _RAND_684 = {1{`RANDOM}};
  rd_D_inBuf_21_validBit = _RAND_684[0:0];
  _RAND_685 = {1{`RANDOM}};
  rd_D_inBuf_21_data = _RAND_685[3:0];
  _RAND_686 = {1{`RANDOM}};
  rd_D_inBuf_22_validBit = _RAND_686[0:0];
  _RAND_687 = {1{`RANDOM}};
  rd_D_inBuf_22_data = _RAND_687[3:0];
  _RAND_688 = {1{`RANDOM}};
  rd_D_inBuf_23_validBit = _RAND_688[0:0];
  _RAND_689 = {1{`RANDOM}};
  rd_D_inBuf_23_data = _RAND_689[3:0];
  _RAND_690 = {1{`RANDOM}};
  rd_D_inBuf_24_validBit = _RAND_690[0:0];
  _RAND_691 = {1{`RANDOM}};
  rd_D_inBuf_24_data = _RAND_691[3:0];
  _RAND_692 = {1{`RANDOM}};
  rd_D_inBuf_25_validBit = _RAND_692[0:0];
  _RAND_693 = {1{`RANDOM}};
  rd_D_inBuf_25_data = _RAND_693[3:0];
  _RAND_694 = {1{`RANDOM}};
  rd_D_inBuf_26_validBit = _RAND_694[0:0];
  _RAND_695 = {1{`RANDOM}};
  rd_D_inBuf_26_data = _RAND_695[3:0];
  _RAND_696 = {1{`RANDOM}};
  rd_D_inBuf_27_validBit = _RAND_696[0:0];
  _RAND_697 = {1{`RANDOM}};
  rd_D_inBuf_27_data = _RAND_697[3:0];
  _RAND_698 = {1{`RANDOM}};
  rd_D_inBuf_28_validBit = _RAND_698[0:0];
  _RAND_699 = {1{`RANDOM}};
  rd_D_inBuf_28_data = _RAND_699[3:0];
  _RAND_700 = {1{`RANDOM}};
  rd_D_inBuf_29_validBit = _RAND_700[0:0];
  _RAND_701 = {1{`RANDOM}};
  rd_D_inBuf_29_data = _RAND_701[3:0];
  _RAND_702 = {1{`RANDOM}};
  rd_D_inBuf_30_validBit = _RAND_702[0:0];
  _RAND_703 = {1{`RANDOM}};
  rd_D_inBuf_30_data = _RAND_703[3:0];
  _RAND_704 = {1{`RANDOM}};
  rd_D_inBuf_31_validBit = _RAND_704[0:0];
  _RAND_705 = {1{`RANDOM}};
  rd_D_inBuf_31_data = _RAND_705[3:0];
  _RAND_706 = {1{`RANDOM}};
  rd_D_inBuf_32_validBit = _RAND_706[0:0];
  _RAND_707 = {1{`RANDOM}};
  rd_D_inBuf_32_data = _RAND_707[3:0];
  _RAND_708 = {1{`RANDOM}};
  rd_D_inBuf_33_validBit = _RAND_708[0:0];
  _RAND_709 = {1{`RANDOM}};
  rd_D_inBuf_33_data = _RAND_709[3:0];
  _RAND_710 = {1{`RANDOM}};
  rd_D_inBuf_34_validBit = _RAND_710[0:0];
  _RAND_711 = {1{`RANDOM}};
  rd_D_inBuf_34_data = _RAND_711[3:0];
  _RAND_712 = {1{`RANDOM}};
  rd_D_inBuf_35_validBit = _RAND_712[0:0];
  _RAND_713 = {1{`RANDOM}};
  rd_D_inBuf_35_data = _RAND_713[3:0];
  _RAND_714 = {1{`RANDOM}};
  rd_D_inBuf_36_validBit = _RAND_714[0:0];
  _RAND_715 = {1{`RANDOM}};
  rd_D_inBuf_36_data = _RAND_715[3:0];
  _RAND_716 = {1{`RANDOM}};
  rd_D_inBuf_37_validBit = _RAND_716[0:0];
  _RAND_717 = {1{`RANDOM}};
  rd_D_inBuf_37_data = _RAND_717[3:0];
  _RAND_718 = {1{`RANDOM}};
  rd_D_inBuf_38_validBit = _RAND_718[0:0];
  _RAND_719 = {1{`RANDOM}};
  rd_D_inBuf_38_data = _RAND_719[3:0];
  _RAND_720 = {1{`RANDOM}};
  rd_D_inBuf_39_validBit = _RAND_720[0:0];
  _RAND_721 = {1{`RANDOM}};
  rd_D_inBuf_39_data = _RAND_721[3:0];
  _RAND_722 = {1{`RANDOM}};
  rd_D_inBuf_40_validBit = _RAND_722[0:0];
  _RAND_723 = {1{`RANDOM}};
  rd_D_inBuf_40_data = _RAND_723[3:0];
  _RAND_724 = {1{`RANDOM}};
  rd_D_inBuf_41_validBit = _RAND_724[0:0];
  _RAND_725 = {1{`RANDOM}};
  rd_D_inBuf_41_data = _RAND_725[3:0];
  _RAND_726 = {1{`RANDOM}};
  rd_D_inBuf_42_validBit = _RAND_726[0:0];
  _RAND_727 = {1{`RANDOM}};
  rd_D_inBuf_42_data = _RAND_727[3:0];
  _RAND_728 = {1{`RANDOM}};
  rd_D_inBuf_43_validBit = _RAND_728[0:0];
  _RAND_729 = {1{`RANDOM}};
  rd_D_inBuf_43_data = _RAND_729[3:0];
  _RAND_730 = {1{`RANDOM}};
  rd_D_inBuf_44_validBit = _RAND_730[0:0];
  _RAND_731 = {1{`RANDOM}};
  rd_D_inBuf_44_data = _RAND_731[3:0];
  _RAND_732 = {1{`RANDOM}};
  rd_D_inBuf_45_validBit = _RAND_732[0:0];
  _RAND_733 = {1{`RANDOM}};
  rd_D_inBuf_45_data = _RAND_733[3:0];
  _RAND_734 = {1{`RANDOM}};
  rd_D_inBuf_46_validBit = _RAND_734[0:0];
  _RAND_735 = {1{`RANDOM}};
  rd_D_inBuf_46_data = _RAND_735[3:0];
  _RAND_736 = {1{`RANDOM}};
  rd_D_inBuf_47_validBit = _RAND_736[0:0];
  _RAND_737 = {1{`RANDOM}};
  rd_D_inBuf_47_data = _RAND_737[3:0];
  _RAND_738 = {1{`RANDOM}};
  rd_D_inBuf_48_validBit = _RAND_738[0:0];
  _RAND_739 = {1{`RANDOM}};
  rd_D_inBuf_48_data = _RAND_739[3:0];
  _RAND_740 = {1{`RANDOM}};
  rd_D_inBuf_49_validBit = _RAND_740[0:0];
  _RAND_741 = {1{`RANDOM}};
  rd_D_inBuf_49_data = _RAND_741[3:0];
  _RAND_742 = {1{`RANDOM}};
  rd_D_inBuf_50_validBit = _RAND_742[0:0];
  _RAND_743 = {1{`RANDOM}};
  rd_D_inBuf_50_data = _RAND_743[3:0];
  _RAND_744 = {1{`RANDOM}};
  rd_D_inBuf_51_validBit = _RAND_744[0:0];
  _RAND_745 = {1{`RANDOM}};
  rd_D_inBuf_51_data = _RAND_745[3:0];
  _RAND_746 = {1{`RANDOM}};
  rd_D_inBuf_52_validBit = _RAND_746[0:0];
  _RAND_747 = {1{`RANDOM}};
  rd_D_inBuf_52_data = _RAND_747[3:0];
  _RAND_748 = {1{`RANDOM}};
  rd_D_inBuf_53_validBit = _RAND_748[0:0];
  _RAND_749 = {1{`RANDOM}};
  rd_D_inBuf_53_data = _RAND_749[3:0];
  _RAND_750 = {1{`RANDOM}};
  rd_D_inBuf_54_validBit = _RAND_750[0:0];
  _RAND_751 = {1{`RANDOM}};
  rd_D_inBuf_54_data = _RAND_751[3:0];
  _RAND_752 = {1{`RANDOM}};
  rd_D_inBuf_55_validBit = _RAND_752[0:0];
  _RAND_753 = {1{`RANDOM}};
  rd_D_inBuf_55_data = _RAND_753[3:0];
  _RAND_754 = {1{`RANDOM}};
  rd_D_inBuf_56_validBit = _RAND_754[0:0];
  _RAND_755 = {1{`RANDOM}};
  rd_D_inBuf_56_data = _RAND_755[3:0];
  _RAND_756 = {1{`RANDOM}};
  rd_D_inBuf_57_validBit = _RAND_756[0:0];
  _RAND_757 = {1{`RANDOM}};
  rd_D_inBuf_57_data = _RAND_757[3:0];
  _RAND_758 = {1{`RANDOM}};
  rd_D_inBuf_58_validBit = _RAND_758[0:0];
  _RAND_759 = {1{`RANDOM}};
  rd_D_inBuf_58_data = _RAND_759[3:0];
  _RAND_760 = {1{`RANDOM}};
  rd_D_inBuf_59_validBit = _RAND_760[0:0];
  _RAND_761 = {1{`RANDOM}};
  rd_D_inBuf_59_data = _RAND_761[3:0];
  _RAND_762 = {1{`RANDOM}};
  rd_D_inBuf_60_validBit = _RAND_762[0:0];
  _RAND_763 = {1{`RANDOM}};
  rd_D_inBuf_60_data = _RAND_763[3:0];
  _RAND_764 = {1{`RANDOM}};
  rd_D_inBuf_61_validBit = _RAND_764[0:0];
  _RAND_765 = {1{`RANDOM}};
  rd_D_inBuf_61_data = _RAND_765[3:0];
  _RAND_766 = {1{`RANDOM}};
  rd_D_inBuf_62_validBit = _RAND_766[0:0];
  _RAND_767 = {1{`RANDOM}};
  rd_D_inBuf_62_data = _RAND_767[3:0];
  _RAND_768 = {1{`RANDOM}};
  rd_D_inBuf_63_validBit = _RAND_768[0:0];
  _RAND_769 = {1{`RANDOM}};
  rd_D_inBuf_63_data = _RAND_769[3:0];
  _RAND_770 = {1{`RANDOM}};
  wr_Addr_outBuf = _RAND_770[7:0];
  _RAND_771 = {1{`RANDOM}};
  wr_D_outBuf_0_validBit = _RAND_771[0:0];
  _RAND_772 = {1{`RANDOM}};
  wr_D_outBuf_0_data = _RAND_772[3:0];
  _RAND_773 = {1{`RANDOM}};
  wr_D_outBuf_1_validBit = _RAND_773[0:0];
  _RAND_774 = {1{`RANDOM}};
  wr_D_outBuf_1_data = _RAND_774[3:0];
  _RAND_775 = {1{`RANDOM}};
  wr_D_outBuf_2_validBit = _RAND_775[0:0];
  _RAND_776 = {1{`RANDOM}};
  wr_D_outBuf_2_data = _RAND_776[3:0];
  _RAND_777 = {1{`RANDOM}};
  wr_D_outBuf_3_validBit = _RAND_777[0:0];
  _RAND_778 = {1{`RANDOM}};
  wr_D_outBuf_3_data = _RAND_778[3:0];
  _RAND_779 = {1{`RANDOM}};
  wr_D_outBuf_4_validBit = _RAND_779[0:0];
  _RAND_780 = {1{`RANDOM}};
  wr_D_outBuf_4_data = _RAND_780[3:0];
  _RAND_781 = {1{`RANDOM}};
  wr_D_outBuf_5_validBit = _RAND_781[0:0];
  _RAND_782 = {1{`RANDOM}};
  wr_D_outBuf_5_data = _RAND_782[3:0];
  _RAND_783 = {1{`RANDOM}};
  wr_D_outBuf_6_validBit = _RAND_783[0:0];
  _RAND_784 = {1{`RANDOM}};
  wr_D_outBuf_6_data = _RAND_784[3:0];
  _RAND_785 = {1{`RANDOM}};
  wr_D_outBuf_7_validBit = _RAND_785[0:0];
  _RAND_786 = {1{`RANDOM}};
  wr_D_outBuf_7_data = _RAND_786[3:0];
  _RAND_787 = {1{`RANDOM}};
  wr_D_outBuf_8_validBit = _RAND_787[0:0];
  _RAND_788 = {1{`RANDOM}};
  wr_D_outBuf_8_data = _RAND_788[3:0];
  _RAND_789 = {1{`RANDOM}};
  wr_D_outBuf_9_validBit = _RAND_789[0:0];
  _RAND_790 = {1{`RANDOM}};
  wr_D_outBuf_9_data = _RAND_790[3:0];
  _RAND_791 = {1{`RANDOM}};
  wr_D_outBuf_10_validBit = _RAND_791[0:0];
  _RAND_792 = {1{`RANDOM}};
  wr_D_outBuf_10_data = _RAND_792[3:0];
  _RAND_793 = {1{`RANDOM}};
  wr_D_outBuf_11_validBit = _RAND_793[0:0];
  _RAND_794 = {1{`RANDOM}};
  wr_D_outBuf_11_data = _RAND_794[3:0];
  _RAND_795 = {1{`RANDOM}};
  wr_D_outBuf_12_validBit = _RAND_795[0:0];
  _RAND_796 = {1{`RANDOM}};
  wr_D_outBuf_12_data = _RAND_796[3:0];
  _RAND_797 = {1{`RANDOM}};
  wr_D_outBuf_13_validBit = _RAND_797[0:0];
  _RAND_798 = {1{`RANDOM}};
  wr_D_outBuf_13_data = _RAND_798[3:0];
  _RAND_799 = {1{`RANDOM}};
  wr_D_outBuf_14_validBit = _RAND_799[0:0];
  _RAND_800 = {1{`RANDOM}};
  wr_D_outBuf_14_data = _RAND_800[3:0];
  _RAND_801 = {1{`RANDOM}};
  wr_D_outBuf_15_validBit = _RAND_801[0:0];
  _RAND_802 = {1{`RANDOM}};
  wr_D_outBuf_15_data = _RAND_802[3:0];
  _RAND_803 = {1{`RANDOM}};
  wr_D_outBuf_16_validBit = _RAND_803[0:0];
  _RAND_804 = {1{`RANDOM}};
  wr_D_outBuf_16_data = _RAND_804[3:0];
  _RAND_805 = {1{`RANDOM}};
  wr_D_outBuf_17_validBit = _RAND_805[0:0];
  _RAND_806 = {1{`RANDOM}};
  wr_D_outBuf_17_data = _RAND_806[3:0];
  _RAND_807 = {1{`RANDOM}};
  wr_D_outBuf_18_validBit = _RAND_807[0:0];
  _RAND_808 = {1{`RANDOM}};
  wr_D_outBuf_18_data = _RAND_808[3:0];
  _RAND_809 = {1{`RANDOM}};
  wr_D_outBuf_19_validBit = _RAND_809[0:0];
  _RAND_810 = {1{`RANDOM}};
  wr_D_outBuf_19_data = _RAND_810[3:0];
  _RAND_811 = {1{`RANDOM}};
  wr_D_outBuf_20_validBit = _RAND_811[0:0];
  _RAND_812 = {1{`RANDOM}};
  wr_D_outBuf_20_data = _RAND_812[3:0];
  _RAND_813 = {1{`RANDOM}};
  wr_D_outBuf_21_validBit = _RAND_813[0:0];
  _RAND_814 = {1{`RANDOM}};
  wr_D_outBuf_21_data = _RAND_814[3:0];
  _RAND_815 = {1{`RANDOM}};
  wr_D_outBuf_22_validBit = _RAND_815[0:0];
  _RAND_816 = {1{`RANDOM}};
  wr_D_outBuf_22_data = _RAND_816[3:0];
  _RAND_817 = {1{`RANDOM}};
  wr_D_outBuf_23_validBit = _RAND_817[0:0];
  _RAND_818 = {1{`RANDOM}};
  wr_D_outBuf_23_data = _RAND_818[3:0];
  _RAND_819 = {1{`RANDOM}};
  wr_D_outBuf_24_validBit = _RAND_819[0:0];
  _RAND_820 = {1{`RANDOM}};
  wr_D_outBuf_24_data = _RAND_820[3:0];
  _RAND_821 = {1{`RANDOM}};
  wr_D_outBuf_25_validBit = _RAND_821[0:0];
  _RAND_822 = {1{`RANDOM}};
  wr_D_outBuf_25_data = _RAND_822[3:0];
  _RAND_823 = {1{`RANDOM}};
  wr_D_outBuf_26_validBit = _RAND_823[0:0];
  _RAND_824 = {1{`RANDOM}};
  wr_D_outBuf_26_data = _RAND_824[3:0];
  _RAND_825 = {1{`RANDOM}};
  wr_D_outBuf_27_validBit = _RAND_825[0:0];
  _RAND_826 = {1{`RANDOM}};
  wr_D_outBuf_27_data = _RAND_826[3:0];
  _RAND_827 = {1{`RANDOM}};
  wr_D_outBuf_28_validBit = _RAND_827[0:0];
  _RAND_828 = {1{`RANDOM}};
  wr_D_outBuf_28_data = _RAND_828[3:0];
  _RAND_829 = {1{`RANDOM}};
  wr_D_outBuf_29_validBit = _RAND_829[0:0];
  _RAND_830 = {1{`RANDOM}};
  wr_D_outBuf_29_data = _RAND_830[3:0];
  _RAND_831 = {1{`RANDOM}};
  wr_D_outBuf_30_validBit = _RAND_831[0:0];
  _RAND_832 = {1{`RANDOM}};
  wr_D_outBuf_30_data = _RAND_832[3:0];
  _RAND_833 = {1{`RANDOM}};
  wr_D_outBuf_31_validBit = _RAND_833[0:0];
  _RAND_834 = {1{`RANDOM}};
  wr_D_outBuf_31_data = _RAND_834[3:0];
  _RAND_835 = {1{`RANDOM}};
  wr_D_outBuf_32_validBit = _RAND_835[0:0];
  _RAND_836 = {1{`RANDOM}};
  wr_D_outBuf_32_data = _RAND_836[3:0];
  _RAND_837 = {1{`RANDOM}};
  wr_D_outBuf_33_validBit = _RAND_837[0:0];
  _RAND_838 = {1{`RANDOM}};
  wr_D_outBuf_33_data = _RAND_838[3:0];
  _RAND_839 = {1{`RANDOM}};
  wr_D_outBuf_34_validBit = _RAND_839[0:0];
  _RAND_840 = {1{`RANDOM}};
  wr_D_outBuf_34_data = _RAND_840[3:0];
  _RAND_841 = {1{`RANDOM}};
  wr_D_outBuf_35_validBit = _RAND_841[0:0];
  _RAND_842 = {1{`RANDOM}};
  wr_D_outBuf_35_data = _RAND_842[3:0];
  _RAND_843 = {1{`RANDOM}};
  wr_D_outBuf_36_validBit = _RAND_843[0:0];
  _RAND_844 = {1{`RANDOM}};
  wr_D_outBuf_36_data = _RAND_844[3:0];
  _RAND_845 = {1{`RANDOM}};
  wr_D_outBuf_37_validBit = _RAND_845[0:0];
  _RAND_846 = {1{`RANDOM}};
  wr_D_outBuf_37_data = _RAND_846[3:0];
  _RAND_847 = {1{`RANDOM}};
  wr_D_outBuf_38_validBit = _RAND_847[0:0];
  _RAND_848 = {1{`RANDOM}};
  wr_D_outBuf_38_data = _RAND_848[3:0];
  _RAND_849 = {1{`RANDOM}};
  wr_D_outBuf_39_validBit = _RAND_849[0:0];
  _RAND_850 = {1{`RANDOM}};
  wr_D_outBuf_39_data = _RAND_850[3:0];
  _RAND_851 = {1{`RANDOM}};
  wr_D_outBuf_40_validBit = _RAND_851[0:0];
  _RAND_852 = {1{`RANDOM}};
  wr_D_outBuf_40_data = _RAND_852[3:0];
  _RAND_853 = {1{`RANDOM}};
  wr_D_outBuf_41_validBit = _RAND_853[0:0];
  _RAND_854 = {1{`RANDOM}};
  wr_D_outBuf_41_data = _RAND_854[3:0];
  _RAND_855 = {1{`RANDOM}};
  wr_D_outBuf_42_validBit = _RAND_855[0:0];
  _RAND_856 = {1{`RANDOM}};
  wr_D_outBuf_42_data = _RAND_856[3:0];
  _RAND_857 = {1{`RANDOM}};
  wr_D_outBuf_43_validBit = _RAND_857[0:0];
  _RAND_858 = {1{`RANDOM}};
  wr_D_outBuf_43_data = _RAND_858[3:0];
  _RAND_859 = {1{`RANDOM}};
  wr_D_outBuf_44_validBit = _RAND_859[0:0];
  _RAND_860 = {1{`RANDOM}};
  wr_D_outBuf_44_data = _RAND_860[3:0];
  _RAND_861 = {1{`RANDOM}};
  wr_D_outBuf_45_validBit = _RAND_861[0:0];
  _RAND_862 = {1{`RANDOM}};
  wr_D_outBuf_45_data = _RAND_862[3:0];
  _RAND_863 = {1{`RANDOM}};
  wr_D_outBuf_46_validBit = _RAND_863[0:0];
  _RAND_864 = {1{`RANDOM}};
  wr_D_outBuf_46_data = _RAND_864[3:0];
  _RAND_865 = {1{`RANDOM}};
  wr_D_outBuf_47_validBit = _RAND_865[0:0];
  _RAND_866 = {1{`RANDOM}};
  wr_D_outBuf_47_data = _RAND_866[3:0];
  _RAND_867 = {1{`RANDOM}};
  wr_D_outBuf_48_validBit = _RAND_867[0:0];
  _RAND_868 = {1{`RANDOM}};
  wr_D_outBuf_48_data = _RAND_868[3:0];
  _RAND_869 = {1{`RANDOM}};
  wr_D_outBuf_49_validBit = _RAND_869[0:0];
  _RAND_870 = {1{`RANDOM}};
  wr_D_outBuf_49_data = _RAND_870[3:0];
  _RAND_871 = {1{`RANDOM}};
  wr_D_outBuf_50_validBit = _RAND_871[0:0];
  _RAND_872 = {1{`RANDOM}};
  wr_D_outBuf_50_data = _RAND_872[3:0];
  _RAND_873 = {1{`RANDOM}};
  wr_D_outBuf_51_validBit = _RAND_873[0:0];
  _RAND_874 = {1{`RANDOM}};
  wr_D_outBuf_51_data = _RAND_874[3:0];
  _RAND_875 = {1{`RANDOM}};
  wr_D_outBuf_52_validBit = _RAND_875[0:0];
  _RAND_876 = {1{`RANDOM}};
  wr_D_outBuf_52_data = _RAND_876[3:0];
  _RAND_877 = {1{`RANDOM}};
  wr_D_outBuf_53_validBit = _RAND_877[0:0];
  _RAND_878 = {1{`RANDOM}};
  wr_D_outBuf_53_data = _RAND_878[3:0];
  _RAND_879 = {1{`RANDOM}};
  wr_D_outBuf_54_validBit = _RAND_879[0:0];
  _RAND_880 = {1{`RANDOM}};
  wr_D_outBuf_54_data = _RAND_880[3:0];
  _RAND_881 = {1{`RANDOM}};
  wr_D_outBuf_55_validBit = _RAND_881[0:0];
  _RAND_882 = {1{`RANDOM}};
  wr_D_outBuf_55_data = _RAND_882[3:0];
  _RAND_883 = {1{`RANDOM}};
  wr_D_outBuf_56_validBit = _RAND_883[0:0];
  _RAND_884 = {1{`RANDOM}};
  wr_D_outBuf_56_data = _RAND_884[3:0];
  _RAND_885 = {1{`RANDOM}};
  wr_D_outBuf_57_validBit = _RAND_885[0:0];
  _RAND_886 = {1{`RANDOM}};
  wr_D_outBuf_57_data = _RAND_886[3:0];
  _RAND_887 = {1{`RANDOM}};
  wr_D_outBuf_58_validBit = _RAND_887[0:0];
  _RAND_888 = {1{`RANDOM}};
  wr_D_outBuf_58_data = _RAND_888[3:0];
  _RAND_889 = {1{`RANDOM}};
  wr_D_outBuf_59_validBit = _RAND_889[0:0];
  _RAND_890 = {1{`RANDOM}};
  wr_D_outBuf_59_data = _RAND_890[3:0];
  _RAND_891 = {1{`RANDOM}};
  wr_D_outBuf_60_validBit = _RAND_891[0:0];
  _RAND_892 = {1{`RANDOM}};
  wr_D_outBuf_60_data = _RAND_892[3:0];
  _RAND_893 = {1{`RANDOM}};
  wr_D_outBuf_61_validBit = _RAND_893[0:0];
  _RAND_894 = {1{`RANDOM}};
  wr_D_outBuf_61_data = _RAND_894[3:0];
  _RAND_895 = {1{`RANDOM}};
  wr_D_outBuf_62_validBit = _RAND_895[0:0];
  _RAND_896 = {1{`RANDOM}};
  wr_D_outBuf_62_data = _RAND_896[3:0];
  _RAND_897 = {1{`RANDOM}};
  wr_D_outBuf_63_validBit = _RAND_897[0:0];
  _RAND_898 = {1{`RANDOM}};
  wr_D_outBuf_63_data = _RAND_898[3:0];
  _RAND_899 = {1{`RANDOM}};
  PCBegin = _RAND_899[7:0];
  _RAND_900 = {1{`RANDOM}};
  AddrBegin = _RAND_900[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
