module CrossBarCell(
  input  [63:0] io_fw_left,
  input  [63:0] io_fw_top,
  output [63:0] io_fw_bottom,
  output [63:0] io_fw_right,
  input         io_sel
);
  assign io_fw_bottom = io_sel ? io_fw_left : io_fw_top; // @[CrossBarSwitchNew.scala 15:17 CrossBarSwitchNew.scala 16:18 CrossBarSwitchNew.scala 18:18]
  assign io_fw_right = io_fw_left; // @[CrossBarSwitchNew.scala 14:15]
endmodule
module CrossBarSwitchNew(
  input         clock,
  input         reset,
  input  [63:0] io_fw_left_0,
  input  [63:0] io_fw_left_1,
  input  [63:0] io_fw_left_2,
  input  [63:0] io_fw_left_3,
  input  [63:0] io_fw_left_4,
  input  [63:0] io_fw_left_5,
  input  [63:0] io_fw_left_6,
  input  [63:0] io_fw_left_7,
  output [63:0] io_fw_bottom_0,
  output [63:0] io_fw_bottom_1,
  output [63:0] io_fw_bottom_2,
  output [63:0] io_fw_bottom_3,
  output [63:0] io_fw_bottom_4,
  output [63:0] io_fw_bottom_5,
  output [63:0] io_fw_bottom_6,
  output [63:0] io_fw_bottom_7,
  input  [2:0]  io_select_0,
  input  [2:0]  io_select_1,
  input  [2:0]  io_select_2,
  input  [2:0]  io_select_3,
  input  [2:0]  io_select_4,
  input  [2:0]  io_select_5,
  input  [2:0]  io_select_6,
  input  [2:0]  io_select_7
);
  wire [63:0] cells_2d_0_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_0_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_0_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_0_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_0_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_1_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_2_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_3_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_4_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_5_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_6_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_7_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_8_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_9_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_10_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_11_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_12_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_13_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_14_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_15_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_16_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_17_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_18_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_19_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_20_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_21_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_22_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_23_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_24_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_25_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_26_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_27_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_28_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_29_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_30_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_31_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_32_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_33_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_34_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_35_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_36_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_37_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_38_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_39_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_40_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_41_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_42_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_43_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_44_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_45_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_46_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_47_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_48_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_49_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_50_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_51_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_52_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_53_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_54_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_55_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_56_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_57_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_58_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_59_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_60_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_61_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_62_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_63_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [7:0] select_onehot_0 = 8'h1 << io_select_0; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_1 = 8'h1 << io_select_1; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_2 = 8'h1 << io_select_2; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_3 = 8'h1 << io_select_3; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_4 = 8'h1 << io_select_4; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_5 = 8'h1 << io_select_5; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_6 = 8'h1 << io_select_6; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_7 = 8'h1 << io_select_7; // @[OneHot.scala 65:12]
  CrossBarCell cells_2d_0 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_0_io_fw_left),
    .io_fw_top(cells_2d_0_io_fw_top),
    .io_fw_bottom(cells_2d_0_io_fw_bottom),
    .io_fw_right(cells_2d_0_io_fw_right),
    .io_sel(cells_2d_0_io_sel)
  );
  CrossBarCell cells_2d_1 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_1_io_fw_left),
    .io_fw_top(cells_2d_1_io_fw_top),
    .io_fw_bottom(cells_2d_1_io_fw_bottom),
    .io_fw_right(cells_2d_1_io_fw_right),
    .io_sel(cells_2d_1_io_sel)
  );
  CrossBarCell cells_2d_2 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_2_io_fw_left),
    .io_fw_top(cells_2d_2_io_fw_top),
    .io_fw_bottom(cells_2d_2_io_fw_bottom),
    .io_fw_right(cells_2d_2_io_fw_right),
    .io_sel(cells_2d_2_io_sel)
  );
  CrossBarCell cells_2d_3 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_3_io_fw_left),
    .io_fw_top(cells_2d_3_io_fw_top),
    .io_fw_bottom(cells_2d_3_io_fw_bottom),
    .io_fw_right(cells_2d_3_io_fw_right),
    .io_sel(cells_2d_3_io_sel)
  );
  CrossBarCell cells_2d_4 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_4_io_fw_left),
    .io_fw_top(cells_2d_4_io_fw_top),
    .io_fw_bottom(cells_2d_4_io_fw_bottom),
    .io_fw_right(cells_2d_4_io_fw_right),
    .io_sel(cells_2d_4_io_sel)
  );
  CrossBarCell cells_2d_5 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_5_io_fw_left),
    .io_fw_top(cells_2d_5_io_fw_top),
    .io_fw_bottom(cells_2d_5_io_fw_bottom),
    .io_fw_right(cells_2d_5_io_fw_right),
    .io_sel(cells_2d_5_io_sel)
  );
  CrossBarCell cells_2d_6 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_6_io_fw_left),
    .io_fw_top(cells_2d_6_io_fw_top),
    .io_fw_bottom(cells_2d_6_io_fw_bottom),
    .io_fw_right(cells_2d_6_io_fw_right),
    .io_sel(cells_2d_6_io_sel)
  );
  CrossBarCell cells_2d_7 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_7_io_fw_left),
    .io_fw_top(cells_2d_7_io_fw_top),
    .io_fw_bottom(cells_2d_7_io_fw_bottom),
    .io_fw_right(cells_2d_7_io_fw_right),
    .io_sel(cells_2d_7_io_sel)
  );
  CrossBarCell cells_2d_8 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_8_io_fw_left),
    .io_fw_top(cells_2d_8_io_fw_top),
    .io_fw_bottom(cells_2d_8_io_fw_bottom),
    .io_fw_right(cells_2d_8_io_fw_right),
    .io_sel(cells_2d_8_io_sel)
  );
  CrossBarCell cells_2d_9 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_9_io_fw_left),
    .io_fw_top(cells_2d_9_io_fw_top),
    .io_fw_bottom(cells_2d_9_io_fw_bottom),
    .io_fw_right(cells_2d_9_io_fw_right),
    .io_sel(cells_2d_9_io_sel)
  );
  CrossBarCell cells_2d_10 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_10_io_fw_left),
    .io_fw_top(cells_2d_10_io_fw_top),
    .io_fw_bottom(cells_2d_10_io_fw_bottom),
    .io_fw_right(cells_2d_10_io_fw_right),
    .io_sel(cells_2d_10_io_sel)
  );
  CrossBarCell cells_2d_11 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_11_io_fw_left),
    .io_fw_top(cells_2d_11_io_fw_top),
    .io_fw_bottom(cells_2d_11_io_fw_bottom),
    .io_fw_right(cells_2d_11_io_fw_right),
    .io_sel(cells_2d_11_io_sel)
  );
  CrossBarCell cells_2d_12 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_12_io_fw_left),
    .io_fw_top(cells_2d_12_io_fw_top),
    .io_fw_bottom(cells_2d_12_io_fw_bottom),
    .io_fw_right(cells_2d_12_io_fw_right),
    .io_sel(cells_2d_12_io_sel)
  );
  CrossBarCell cells_2d_13 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_13_io_fw_left),
    .io_fw_top(cells_2d_13_io_fw_top),
    .io_fw_bottom(cells_2d_13_io_fw_bottom),
    .io_fw_right(cells_2d_13_io_fw_right),
    .io_sel(cells_2d_13_io_sel)
  );
  CrossBarCell cells_2d_14 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_14_io_fw_left),
    .io_fw_top(cells_2d_14_io_fw_top),
    .io_fw_bottom(cells_2d_14_io_fw_bottom),
    .io_fw_right(cells_2d_14_io_fw_right),
    .io_sel(cells_2d_14_io_sel)
  );
  CrossBarCell cells_2d_15 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_15_io_fw_left),
    .io_fw_top(cells_2d_15_io_fw_top),
    .io_fw_bottom(cells_2d_15_io_fw_bottom),
    .io_fw_right(cells_2d_15_io_fw_right),
    .io_sel(cells_2d_15_io_sel)
  );
  CrossBarCell cells_2d_16 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_16_io_fw_left),
    .io_fw_top(cells_2d_16_io_fw_top),
    .io_fw_bottom(cells_2d_16_io_fw_bottom),
    .io_fw_right(cells_2d_16_io_fw_right),
    .io_sel(cells_2d_16_io_sel)
  );
  CrossBarCell cells_2d_17 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_17_io_fw_left),
    .io_fw_top(cells_2d_17_io_fw_top),
    .io_fw_bottom(cells_2d_17_io_fw_bottom),
    .io_fw_right(cells_2d_17_io_fw_right),
    .io_sel(cells_2d_17_io_sel)
  );
  CrossBarCell cells_2d_18 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_18_io_fw_left),
    .io_fw_top(cells_2d_18_io_fw_top),
    .io_fw_bottom(cells_2d_18_io_fw_bottom),
    .io_fw_right(cells_2d_18_io_fw_right),
    .io_sel(cells_2d_18_io_sel)
  );
  CrossBarCell cells_2d_19 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_19_io_fw_left),
    .io_fw_top(cells_2d_19_io_fw_top),
    .io_fw_bottom(cells_2d_19_io_fw_bottom),
    .io_fw_right(cells_2d_19_io_fw_right),
    .io_sel(cells_2d_19_io_sel)
  );
  CrossBarCell cells_2d_20 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_20_io_fw_left),
    .io_fw_top(cells_2d_20_io_fw_top),
    .io_fw_bottom(cells_2d_20_io_fw_bottom),
    .io_fw_right(cells_2d_20_io_fw_right),
    .io_sel(cells_2d_20_io_sel)
  );
  CrossBarCell cells_2d_21 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_21_io_fw_left),
    .io_fw_top(cells_2d_21_io_fw_top),
    .io_fw_bottom(cells_2d_21_io_fw_bottom),
    .io_fw_right(cells_2d_21_io_fw_right),
    .io_sel(cells_2d_21_io_sel)
  );
  CrossBarCell cells_2d_22 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_22_io_fw_left),
    .io_fw_top(cells_2d_22_io_fw_top),
    .io_fw_bottom(cells_2d_22_io_fw_bottom),
    .io_fw_right(cells_2d_22_io_fw_right),
    .io_sel(cells_2d_22_io_sel)
  );
  CrossBarCell cells_2d_23 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_23_io_fw_left),
    .io_fw_top(cells_2d_23_io_fw_top),
    .io_fw_bottom(cells_2d_23_io_fw_bottom),
    .io_fw_right(cells_2d_23_io_fw_right),
    .io_sel(cells_2d_23_io_sel)
  );
  CrossBarCell cells_2d_24 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_24_io_fw_left),
    .io_fw_top(cells_2d_24_io_fw_top),
    .io_fw_bottom(cells_2d_24_io_fw_bottom),
    .io_fw_right(cells_2d_24_io_fw_right),
    .io_sel(cells_2d_24_io_sel)
  );
  CrossBarCell cells_2d_25 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_25_io_fw_left),
    .io_fw_top(cells_2d_25_io_fw_top),
    .io_fw_bottom(cells_2d_25_io_fw_bottom),
    .io_fw_right(cells_2d_25_io_fw_right),
    .io_sel(cells_2d_25_io_sel)
  );
  CrossBarCell cells_2d_26 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_26_io_fw_left),
    .io_fw_top(cells_2d_26_io_fw_top),
    .io_fw_bottom(cells_2d_26_io_fw_bottom),
    .io_fw_right(cells_2d_26_io_fw_right),
    .io_sel(cells_2d_26_io_sel)
  );
  CrossBarCell cells_2d_27 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_27_io_fw_left),
    .io_fw_top(cells_2d_27_io_fw_top),
    .io_fw_bottom(cells_2d_27_io_fw_bottom),
    .io_fw_right(cells_2d_27_io_fw_right),
    .io_sel(cells_2d_27_io_sel)
  );
  CrossBarCell cells_2d_28 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_28_io_fw_left),
    .io_fw_top(cells_2d_28_io_fw_top),
    .io_fw_bottom(cells_2d_28_io_fw_bottom),
    .io_fw_right(cells_2d_28_io_fw_right),
    .io_sel(cells_2d_28_io_sel)
  );
  CrossBarCell cells_2d_29 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_29_io_fw_left),
    .io_fw_top(cells_2d_29_io_fw_top),
    .io_fw_bottom(cells_2d_29_io_fw_bottom),
    .io_fw_right(cells_2d_29_io_fw_right),
    .io_sel(cells_2d_29_io_sel)
  );
  CrossBarCell cells_2d_30 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_30_io_fw_left),
    .io_fw_top(cells_2d_30_io_fw_top),
    .io_fw_bottom(cells_2d_30_io_fw_bottom),
    .io_fw_right(cells_2d_30_io_fw_right),
    .io_sel(cells_2d_30_io_sel)
  );
  CrossBarCell cells_2d_31 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_31_io_fw_left),
    .io_fw_top(cells_2d_31_io_fw_top),
    .io_fw_bottom(cells_2d_31_io_fw_bottom),
    .io_fw_right(cells_2d_31_io_fw_right),
    .io_sel(cells_2d_31_io_sel)
  );
  CrossBarCell cells_2d_32 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_32_io_fw_left),
    .io_fw_top(cells_2d_32_io_fw_top),
    .io_fw_bottom(cells_2d_32_io_fw_bottom),
    .io_fw_right(cells_2d_32_io_fw_right),
    .io_sel(cells_2d_32_io_sel)
  );
  CrossBarCell cells_2d_33 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_33_io_fw_left),
    .io_fw_top(cells_2d_33_io_fw_top),
    .io_fw_bottom(cells_2d_33_io_fw_bottom),
    .io_fw_right(cells_2d_33_io_fw_right),
    .io_sel(cells_2d_33_io_sel)
  );
  CrossBarCell cells_2d_34 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_34_io_fw_left),
    .io_fw_top(cells_2d_34_io_fw_top),
    .io_fw_bottom(cells_2d_34_io_fw_bottom),
    .io_fw_right(cells_2d_34_io_fw_right),
    .io_sel(cells_2d_34_io_sel)
  );
  CrossBarCell cells_2d_35 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_35_io_fw_left),
    .io_fw_top(cells_2d_35_io_fw_top),
    .io_fw_bottom(cells_2d_35_io_fw_bottom),
    .io_fw_right(cells_2d_35_io_fw_right),
    .io_sel(cells_2d_35_io_sel)
  );
  CrossBarCell cells_2d_36 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_36_io_fw_left),
    .io_fw_top(cells_2d_36_io_fw_top),
    .io_fw_bottom(cells_2d_36_io_fw_bottom),
    .io_fw_right(cells_2d_36_io_fw_right),
    .io_sel(cells_2d_36_io_sel)
  );
  CrossBarCell cells_2d_37 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_37_io_fw_left),
    .io_fw_top(cells_2d_37_io_fw_top),
    .io_fw_bottom(cells_2d_37_io_fw_bottom),
    .io_fw_right(cells_2d_37_io_fw_right),
    .io_sel(cells_2d_37_io_sel)
  );
  CrossBarCell cells_2d_38 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_38_io_fw_left),
    .io_fw_top(cells_2d_38_io_fw_top),
    .io_fw_bottom(cells_2d_38_io_fw_bottom),
    .io_fw_right(cells_2d_38_io_fw_right),
    .io_sel(cells_2d_38_io_sel)
  );
  CrossBarCell cells_2d_39 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_39_io_fw_left),
    .io_fw_top(cells_2d_39_io_fw_top),
    .io_fw_bottom(cells_2d_39_io_fw_bottom),
    .io_fw_right(cells_2d_39_io_fw_right),
    .io_sel(cells_2d_39_io_sel)
  );
  CrossBarCell cells_2d_40 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_40_io_fw_left),
    .io_fw_top(cells_2d_40_io_fw_top),
    .io_fw_bottom(cells_2d_40_io_fw_bottom),
    .io_fw_right(cells_2d_40_io_fw_right),
    .io_sel(cells_2d_40_io_sel)
  );
  CrossBarCell cells_2d_41 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_41_io_fw_left),
    .io_fw_top(cells_2d_41_io_fw_top),
    .io_fw_bottom(cells_2d_41_io_fw_bottom),
    .io_fw_right(cells_2d_41_io_fw_right),
    .io_sel(cells_2d_41_io_sel)
  );
  CrossBarCell cells_2d_42 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_42_io_fw_left),
    .io_fw_top(cells_2d_42_io_fw_top),
    .io_fw_bottom(cells_2d_42_io_fw_bottom),
    .io_fw_right(cells_2d_42_io_fw_right),
    .io_sel(cells_2d_42_io_sel)
  );
  CrossBarCell cells_2d_43 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_43_io_fw_left),
    .io_fw_top(cells_2d_43_io_fw_top),
    .io_fw_bottom(cells_2d_43_io_fw_bottom),
    .io_fw_right(cells_2d_43_io_fw_right),
    .io_sel(cells_2d_43_io_sel)
  );
  CrossBarCell cells_2d_44 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_44_io_fw_left),
    .io_fw_top(cells_2d_44_io_fw_top),
    .io_fw_bottom(cells_2d_44_io_fw_bottom),
    .io_fw_right(cells_2d_44_io_fw_right),
    .io_sel(cells_2d_44_io_sel)
  );
  CrossBarCell cells_2d_45 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_45_io_fw_left),
    .io_fw_top(cells_2d_45_io_fw_top),
    .io_fw_bottom(cells_2d_45_io_fw_bottom),
    .io_fw_right(cells_2d_45_io_fw_right),
    .io_sel(cells_2d_45_io_sel)
  );
  CrossBarCell cells_2d_46 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_46_io_fw_left),
    .io_fw_top(cells_2d_46_io_fw_top),
    .io_fw_bottom(cells_2d_46_io_fw_bottom),
    .io_fw_right(cells_2d_46_io_fw_right),
    .io_sel(cells_2d_46_io_sel)
  );
  CrossBarCell cells_2d_47 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_47_io_fw_left),
    .io_fw_top(cells_2d_47_io_fw_top),
    .io_fw_bottom(cells_2d_47_io_fw_bottom),
    .io_fw_right(cells_2d_47_io_fw_right),
    .io_sel(cells_2d_47_io_sel)
  );
  CrossBarCell cells_2d_48 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_48_io_fw_left),
    .io_fw_top(cells_2d_48_io_fw_top),
    .io_fw_bottom(cells_2d_48_io_fw_bottom),
    .io_fw_right(cells_2d_48_io_fw_right),
    .io_sel(cells_2d_48_io_sel)
  );
  CrossBarCell cells_2d_49 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_49_io_fw_left),
    .io_fw_top(cells_2d_49_io_fw_top),
    .io_fw_bottom(cells_2d_49_io_fw_bottom),
    .io_fw_right(cells_2d_49_io_fw_right),
    .io_sel(cells_2d_49_io_sel)
  );
  CrossBarCell cells_2d_50 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_50_io_fw_left),
    .io_fw_top(cells_2d_50_io_fw_top),
    .io_fw_bottom(cells_2d_50_io_fw_bottom),
    .io_fw_right(cells_2d_50_io_fw_right),
    .io_sel(cells_2d_50_io_sel)
  );
  CrossBarCell cells_2d_51 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_51_io_fw_left),
    .io_fw_top(cells_2d_51_io_fw_top),
    .io_fw_bottom(cells_2d_51_io_fw_bottom),
    .io_fw_right(cells_2d_51_io_fw_right),
    .io_sel(cells_2d_51_io_sel)
  );
  CrossBarCell cells_2d_52 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_52_io_fw_left),
    .io_fw_top(cells_2d_52_io_fw_top),
    .io_fw_bottom(cells_2d_52_io_fw_bottom),
    .io_fw_right(cells_2d_52_io_fw_right),
    .io_sel(cells_2d_52_io_sel)
  );
  CrossBarCell cells_2d_53 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_53_io_fw_left),
    .io_fw_top(cells_2d_53_io_fw_top),
    .io_fw_bottom(cells_2d_53_io_fw_bottom),
    .io_fw_right(cells_2d_53_io_fw_right),
    .io_sel(cells_2d_53_io_sel)
  );
  CrossBarCell cells_2d_54 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_54_io_fw_left),
    .io_fw_top(cells_2d_54_io_fw_top),
    .io_fw_bottom(cells_2d_54_io_fw_bottom),
    .io_fw_right(cells_2d_54_io_fw_right),
    .io_sel(cells_2d_54_io_sel)
  );
  CrossBarCell cells_2d_55 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_55_io_fw_left),
    .io_fw_top(cells_2d_55_io_fw_top),
    .io_fw_bottom(cells_2d_55_io_fw_bottom),
    .io_fw_right(cells_2d_55_io_fw_right),
    .io_sel(cells_2d_55_io_sel)
  );
  CrossBarCell cells_2d_56 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_56_io_fw_left),
    .io_fw_top(cells_2d_56_io_fw_top),
    .io_fw_bottom(cells_2d_56_io_fw_bottom),
    .io_fw_right(cells_2d_56_io_fw_right),
    .io_sel(cells_2d_56_io_sel)
  );
  CrossBarCell cells_2d_57 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_57_io_fw_left),
    .io_fw_top(cells_2d_57_io_fw_top),
    .io_fw_bottom(cells_2d_57_io_fw_bottom),
    .io_fw_right(cells_2d_57_io_fw_right),
    .io_sel(cells_2d_57_io_sel)
  );
  CrossBarCell cells_2d_58 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_58_io_fw_left),
    .io_fw_top(cells_2d_58_io_fw_top),
    .io_fw_bottom(cells_2d_58_io_fw_bottom),
    .io_fw_right(cells_2d_58_io_fw_right),
    .io_sel(cells_2d_58_io_sel)
  );
  CrossBarCell cells_2d_59 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_59_io_fw_left),
    .io_fw_top(cells_2d_59_io_fw_top),
    .io_fw_bottom(cells_2d_59_io_fw_bottom),
    .io_fw_right(cells_2d_59_io_fw_right),
    .io_sel(cells_2d_59_io_sel)
  );
  CrossBarCell cells_2d_60 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_60_io_fw_left),
    .io_fw_top(cells_2d_60_io_fw_top),
    .io_fw_bottom(cells_2d_60_io_fw_bottom),
    .io_fw_right(cells_2d_60_io_fw_right),
    .io_sel(cells_2d_60_io_sel)
  );
  CrossBarCell cells_2d_61 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_61_io_fw_left),
    .io_fw_top(cells_2d_61_io_fw_top),
    .io_fw_bottom(cells_2d_61_io_fw_bottom),
    .io_fw_right(cells_2d_61_io_fw_right),
    .io_sel(cells_2d_61_io_sel)
  );
  CrossBarCell cells_2d_62 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_62_io_fw_left),
    .io_fw_top(cells_2d_62_io_fw_top),
    .io_fw_bottom(cells_2d_62_io_fw_bottom),
    .io_fw_right(cells_2d_62_io_fw_right),
    .io_sel(cells_2d_62_io_sel)
  );
  CrossBarCell cells_2d_63 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_63_io_fw_left),
    .io_fw_top(cells_2d_63_io_fw_top),
    .io_fw_bottom(cells_2d_63_io_fw_bottom),
    .io_fw_right(cells_2d_63_io_fw_right),
    .io_sel(cells_2d_63_io_sel)
  );
  assign io_fw_bottom_0 = cells_2d_56_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_1 = cells_2d_57_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_2 = cells_2d_58_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_3 = cells_2d_59_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_4 = cells_2d_60_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_5 = cells_2d_61_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_6 = cells_2d_62_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_7 = cells_2d_63_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign cells_2d_0_io_fw_left = io_fw_left_0; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_0_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_0_io_sel = select_onehot_0[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_1_io_fw_left = cells_2d_0_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_1_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_1_io_sel = select_onehot_1[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_2_io_fw_left = cells_2d_1_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_2_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_2_io_sel = select_onehot_2[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_3_io_fw_left = cells_2d_2_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_3_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_3_io_sel = select_onehot_3[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_4_io_fw_left = cells_2d_3_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_4_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_4_io_sel = select_onehot_4[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_5_io_fw_left = cells_2d_4_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_5_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_5_io_sel = select_onehot_5[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_6_io_fw_left = cells_2d_5_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_6_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_6_io_sel = select_onehot_6[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_7_io_fw_left = cells_2d_6_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_7_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_7_io_sel = select_onehot_7[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_8_io_fw_left = io_fw_left_1; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_8_io_fw_top = cells_2d_0_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_8_io_sel = select_onehot_0[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_9_io_fw_left = cells_2d_8_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_9_io_fw_top = cells_2d_1_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_9_io_sel = select_onehot_1[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_10_io_fw_left = cells_2d_9_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_10_io_fw_top = cells_2d_2_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_10_io_sel = select_onehot_2[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_11_io_fw_left = cells_2d_10_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_11_io_fw_top = cells_2d_3_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_11_io_sel = select_onehot_3[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_12_io_fw_left = cells_2d_11_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_12_io_fw_top = cells_2d_4_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_12_io_sel = select_onehot_4[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_13_io_fw_left = cells_2d_12_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_13_io_fw_top = cells_2d_5_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_13_io_sel = select_onehot_5[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_14_io_fw_left = cells_2d_13_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_14_io_fw_top = cells_2d_6_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_14_io_sel = select_onehot_6[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_15_io_fw_left = cells_2d_14_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_15_io_fw_top = cells_2d_7_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_15_io_sel = select_onehot_7[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_16_io_fw_left = io_fw_left_2; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_16_io_fw_top = cells_2d_8_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_16_io_sel = select_onehot_0[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_17_io_fw_left = cells_2d_16_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_17_io_fw_top = cells_2d_9_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_17_io_sel = select_onehot_1[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_18_io_fw_left = cells_2d_17_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_18_io_fw_top = cells_2d_10_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_18_io_sel = select_onehot_2[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_19_io_fw_left = cells_2d_18_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_19_io_fw_top = cells_2d_11_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_19_io_sel = select_onehot_3[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_20_io_fw_left = cells_2d_19_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_20_io_fw_top = cells_2d_12_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_20_io_sel = select_onehot_4[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_21_io_fw_left = cells_2d_20_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_21_io_fw_top = cells_2d_13_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_21_io_sel = select_onehot_5[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_22_io_fw_left = cells_2d_21_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_22_io_fw_top = cells_2d_14_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_22_io_sel = select_onehot_6[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_23_io_fw_left = cells_2d_22_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_23_io_fw_top = cells_2d_15_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_23_io_sel = select_onehot_7[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_24_io_fw_left = io_fw_left_3; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_24_io_fw_top = cells_2d_16_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_24_io_sel = select_onehot_0[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_25_io_fw_left = cells_2d_24_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_25_io_fw_top = cells_2d_17_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_25_io_sel = select_onehot_1[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_26_io_fw_left = cells_2d_25_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_26_io_fw_top = cells_2d_18_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_26_io_sel = select_onehot_2[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_27_io_fw_left = cells_2d_26_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_27_io_fw_top = cells_2d_19_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_27_io_sel = select_onehot_3[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_28_io_fw_left = cells_2d_27_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_28_io_fw_top = cells_2d_20_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_28_io_sel = select_onehot_4[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_29_io_fw_left = cells_2d_28_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_29_io_fw_top = cells_2d_21_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_29_io_sel = select_onehot_5[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_30_io_fw_left = cells_2d_29_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_30_io_fw_top = cells_2d_22_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_30_io_sel = select_onehot_6[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_31_io_fw_left = cells_2d_30_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_31_io_fw_top = cells_2d_23_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_31_io_sel = select_onehot_7[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_32_io_fw_left = io_fw_left_4; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_32_io_fw_top = cells_2d_24_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_32_io_sel = select_onehot_0[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_33_io_fw_left = cells_2d_32_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_33_io_fw_top = cells_2d_25_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_33_io_sel = select_onehot_1[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_34_io_fw_left = cells_2d_33_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_34_io_fw_top = cells_2d_26_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_34_io_sel = select_onehot_2[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_35_io_fw_left = cells_2d_34_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_35_io_fw_top = cells_2d_27_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_35_io_sel = select_onehot_3[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_36_io_fw_left = cells_2d_35_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_36_io_fw_top = cells_2d_28_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_36_io_sel = select_onehot_4[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_37_io_fw_left = cells_2d_36_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_37_io_fw_top = cells_2d_29_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_37_io_sel = select_onehot_5[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_38_io_fw_left = cells_2d_37_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_38_io_fw_top = cells_2d_30_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_38_io_sel = select_onehot_6[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_39_io_fw_left = cells_2d_38_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_39_io_fw_top = cells_2d_31_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_39_io_sel = select_onehot_7[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_40_io_fw_left = io_fw_left_5; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_40_io_fw_top = cells_2d_32_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_40_io_sel = select_onehot_0[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_41_io_fw_left = cells_2d_40_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_41_io_fw_top = cells_2d_33_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_41_io_sel = select_onehot_1[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_42_io_fw_left = cells_2d_41_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_42_io_fw_top = cells_2d_34_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_42_io_sel = select_onehot_2[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_43_io_fw_left = cells_2d_42_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_43_io_fw_top = cells_2d_35_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_43_io_sel = select_onehot_3[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_44_io_fw_left = cells_2d_43_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_44_io_fw_top = cells_2d_36_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_44_io_sel = select_onehot_4[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_45_io_fw_left = cells_2d_44_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_45_io_fw_top = cells_2d_37_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_45_io_sel = select_onehot_5[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_46_io_fw_left = cells_2d_45_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_46_io_fw_top = cells_2d_38_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_46_io_sel = select_onehot_6[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_47_io_fw_left = cells_2d_46_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_47_io_fw_top = cells_2d_39_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_47_io_sel = select_onehot_7[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_48_io_fw_left = io_fw_left_6; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_48_io_fw_top = cells_2d_40_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_48_io_sel = select_onehot_0[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_49_io_fw_left = cells_2d_48_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_49_io_fw_top = cells_2d_41_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_49_io_sel = select_onehot_1[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_50_io_fw_left = cells_2d_49_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_50_io_fw_top = cells_2d_42_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_50_io_sel = select_onehot_2[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_51_io_fw_left = cells_2d_50_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_51_io_fw_top = cells_2d_43_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_51_io_sel = select_onehot_3[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_52_io_fw_left = cells_2d_51_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_52_io_fw_top = cells_2d_44_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_52_io_sel = select_onehot_4[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_53_io_fw_left = cells_2d_52_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_53_io_fw_top = cells_2d_45_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_53_io_sel = select_onehot_5[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_54_io_fw_left = cells_2d_53_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_54_io_fw_top = cells_2d_46_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_54_io_sel = select_onehot_6[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_55_io_fw_left = cells_2d_54_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_55_io_fw_top = cells_2d_47_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_55_io_sel = select_onehot_7[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_56_io_fw_left = io_fw_left_7; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_56_io_fw_top = cells_2d_48_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_56_io_sel = select_onehot_0[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_57_io_fw_left = cells_2d_56_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_57_io_fw_top = cells_2d_49_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_57_io_sel = select_onehot_1[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_58_io_fw_left = cells_2d_57_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_58_io_fw_top = cells_2d_50_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_58_io_sel = select_onehot_2[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_59_io_fw_left = cells_2d_58_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_59_io_fw_top = cells_2d_51_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_59_io_sel = select_onehot_3[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_60_io_fw_left = cells_2d_59_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_60_io_fw_top = cells_2d_52_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_60_io_sel = select_onehot_4[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_61_io_fw_left = cells_2d_60_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_61_io_fw_top = cells_2d_53_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_61_io_sel = select_onehot_5[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_62_io_fw_left = cells_2d_61_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_62_io_fw_top = cells_2d_54_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_62_io_sel = select_onehot_6[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_63_io_fw_left = cells_2d_62_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_63_io_fw_top = cells_2d_55_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_63_io_sel = select_onehot_7[7]; // @[CrossBarSwitchNew.scala 70:44]
endmodule
