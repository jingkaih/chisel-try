module CrossBarCell(
  input  [63:0] io_fw_left,
  input  [63:0] io_fw_top,
  output [63:0] io_fw_bottom,
  output [63:0] io_fw_right,
  input         io_sel
);
  assign io_fw_bottom = io_sel ? io_fw_left : io_fw_top; // @[CrossBarSwitchNew.scala 15:17 CrossBarSwitchNew.scala 16:18 CrossBarSwitchNew.scala 18:18]
  assign io_fw_right = io_fw_left; // @[CrossBarSwitchNew.scala 14:15]
endmodule
module CrossBarSwitchNew(
  input  [63:0] io_fw_left_0,
  input  [63:0] io_fw_left_1,
  input  [63:0] io_fw_left_2,
  input  [63:0] io_fw_left_3,
  input  [63:0] io_fw_left_4,
  input  [63:0] io_fw_left_5,
  input  [63:0] io_fw_left_6,
  input  [63:0] io_fw_left_7,
  output [63:0] io_fw_bottom_0,
  output [63:0] io_fw_bottom_1,
  output [63:0] io_fw_bottom_2,
  output [63:0] io_fw_bottom_3,
  output [63:0] io_fw_bottom_4,
  output [63:0] io_fw_bottom_5,
  output [63:0] io_fw_bottom_6,
  output [63:0] io_fw_bottom_7,
  input  [2:0]  io_select_0,
  input  [2:0]  io_select_1,
  input  [2:0]  io_select_2,
  input  [2:0]  io_select_3,
  input  [2:0]  io_select_4,
  input  [2:0]  io_select_5,
  input  [2:0]  io_select_6,
  input  [2:0]  io_select_7
);
  wire [63:0] cells_2d_0_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_0_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_0_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_0_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_0_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_1_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_1_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_2_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_2_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_3_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_3_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_4_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_4_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_5_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_5_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_6_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_6_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_7_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_7_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_8_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_8_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_9_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_9_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_10_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_10_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_11_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_11_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_12_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_12_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_13_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_13_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_14_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_14_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_15_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_15_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_16_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_16_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_17_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_17_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_18_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_18_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_19_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_19_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_20_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_20_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_21_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_21_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_22_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_22_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_23_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_23_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_24_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_24_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_25_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_25_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_26_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_26_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_27_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_27_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_28_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_28_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_29_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_29_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_30_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_30_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_31_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_31_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_32_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_32_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_33_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_33_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_34_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_34_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_35_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_35_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_36_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_36_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_37_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_37_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_38_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_38_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_39_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_39_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_40_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_40_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_41_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_41_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_42_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_42_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_43_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_43_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_44_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_44_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_45_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_45_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_46_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_46_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_47_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_47_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_48_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_48_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_49_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_49_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_50_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_50_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_51_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_51_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_52_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_52_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_53_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_53_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_54_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_54_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_55_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_55_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_56_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_56_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_57_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_57_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_58_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_58_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_59_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_59_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_60_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_60_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_61_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_61_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_62_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_62_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_left; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_top; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_bottom; // @[CrossBarSwitchNew.scala 38:53]
  wire [63:0] cells_2d_63_io_fw_right; // @[CrossBarSwitchNew.scala 38:53]
  wire  cells_2d_63_io_sel; // @[CrossBarSwitchNew.scala 38:53]
  wire [7:0] select_onehot_0 = 8'h1 << io_select_0; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_1 = 8'h1 << io_select_1; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_2 = 8'h1 << io_select_2; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_3 = 8'h1 << io_select_3; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_4 = 8'h1 << io_select_4; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_5 = 8'h1 << io_select_5; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_6 = 8'h1 << io_select_6; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_7 = 8'h1 << io_select_7; // @[OneHot.scala 65:12]
  CrossBarCell cells_2d_0 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_0_io_fw_left),
    .io_fw_top(cells_2d_0_io_fw_top),
    .io_fw_bottom(cells_2d_0_io_fw_bottom),
    .io_fw_right(cells_2d_0_io_fw_right),
    .io_sel(cells_2d_0_io_sel)
  );
  CrossBarCell cells_2d_1 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_1_io_fw_left),
    .io_fw_top(cells_2d_1_io_fw_top),
    .io_fw_bottom(cells_2d_1_io_fw_bottom),
    .io_fw_right(cells_2d_1_io_fw_right),
    .io_sel(cells_2d_1_io_sel)
  );
  CrossBarCell cells_2d_2 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_2_io_fw_left),
    .io_fw_top(cells_2d_2_io_fw_top),
    .io_fw_bottom(cells_2d_2_io_fw_bottom),
    .io_fw_right(cells_2d_2_io_fw_right),
    .io_sel(cells_2d_2_io_sel)
  );
  CrossBarCell cells_2d_3 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_3_io_fw_left),
    .io_fw_top(cells_2d_3_io_fw_top),
    .io_fw_bottom(cells_2d_3_io_fw_bottom),
    .io_fw_right(cells_2d_3_io_fw_right),
    .io_sel(cells_2d_3_io_sel)
  );
  CrossBarCell cells_2d_4 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_4_io_fw_left),
    .io_fw_top(cells_2d_4_io_fw_top),
    .io_fw_bottom(cells_2d_4_io_fw_bottom),
    .io_fw_right(cells_2d_4_io_fw_right),
    .io_sel(cells_2d_4_io_sel)
  );
  CrossBarCell cells_2d_5 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_5_io_fw_left),
    .io_fw_top(cells_2d_5_io_fw_top),
    .io_fw_bottom(cells_2d_5_io_fw_bottom),
    .io_fw_right(cells_2d_5_io_fw_right),
    .io_sel(cells_2d_5_io_sel)
  );
  CrossBarCell cells_2d_6 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_6_io_fw_left),
    .io_fw_top(cells_2d_6_io_fw_top),
    .io_fw_bottom(cells_2d_6_io_fw_bottom),
    .io_fw_right(cells_2d_6_io_fw_right),
    .io_sel(cells_2d_6_io_sel)
  );
  CrossBarCell cells_2d_7 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_7_io_fw_left),
    .io_fw_top(cells_2d_7_io_fw_top),
    .io_fw_bottom(cells_2d_7_io_fw_bottom),
    .io_fw_right(cells_2d_7_io_fw_right),
    .io_sel(cells_2d_7_io_sel)
  );
  CrossBarCell cells_2d_8 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_8_io_fw_left),
    .io_fw_top(cells_2d_8_io_fw_top),
    .io_fw_bottom(cells_2d_8_io_fw_bottom),
    .io_fw_right(cells_2d_8_io_fw_right),
    .io_sel(cells_2d_8_io_sel)
  );
  CrossBarCell cells_2d_9 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_9_io_fw_left),
    .io_fw_top(cells_2d_9_io_fw_top),
    .io_fw_bottom(cells_2d_9_io_fw_bottom),
    .io_fw_right(cells_2d_9_io_fw_right),
    .io_sel(cells_2d_9_io_sel)
  );
  CrossBarCell cells_2d_10 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_10_io_fw_left),
    .io_fw_top(cells_2d_10_io_fw_top),
    .io_fw_bottom(cells_2d_10_io_fw_bottom),
    .io_fw_right(cells_2d_10_io_fw_right),
    .io_sel(cells_2d_10_io_sel)
  );
  CrossBarCell cells_2d_11 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_11_io_fw_left),
    .io_fw_top(cells_2d_11_io_fw_top),
    .io_fw_bottom(cells_2d_11_io_fw_bottom),
    .io_fw_right(cells_2d_11_io_fw_right),
    .io_sel(cells_2d_11_io_sel)
  );
  CrossBarCell cells_2d_12 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_12_io_fw_left),
    .io_fw_top(cells_2d_12_io_fw_top),
    .io_fw_bottom(cells_2d_12_io_fw_bottom),
    .io_fw_right(cells_2d_12_io_fw_right),
    .io_sel(cells_2d_12_io_sel)
  );
  CrossBarCell cells_2d_13 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_13_io_fw_left),
    .io_fw_top(cells_2d_13_io_fw_top),
    .io_fw_bottom(cells_2d_13_io_fw_bottom),
    .io_fw_right(cells_2d_13_io_fw_right),
    .io_sel(cells_2d_13_io_sel)
  );
  CrossBarCell cells_2d_14 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_14_io_fw_left),
    .io_fw_top(cells_2d_14_io_fw_top),
    .io_fw_bottom(cells_2d_14_io_fw_bottom),
    .io_fw_right(cells_2d_14_io_fw_right),
    .io_sel(cells_2d_14_io_sel)
  );
  CrossBarCell cells_2d_15 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_15_io_fw_left),
    .io_fw_top(cells_2d_15_io_fw_top),
    .io_fw_bottom(cells_2d_15_io_fw_bottom),
    .io_fw_right(cells_2d_15_io_fw_right),
    .io_sel(cells_2d_15_io_sel)
  );
  CrossBarCell cells_2d_16 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_16_io_fw_left),
    .io_fw_top(cells_2d_16_io_fw_top),
    .io_fw_bottom(cells_2d_16_io_fw_bottom),
    .io_fw_right(cells_2d_16_io_fw_right),
    .io_sel(cells_2d_16_io_sel)
  );
  CrossBarCell cells_2d_17 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_17_io_fw_left),
    .io_fw_top(cells_2d_17_io_fw_top),
    .io_fw_bottom(cells_2d_17_io_fw_bottom),
    .io_fw_right(cells_2d_17_io_fw_right),
    .io_sel(cells_2d_17_io_sel)
  );
  CrossBarCell cells_2d_18 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_18_io_fw_left),
    .io_fw_top(cells_2d_18_io_fw_top),
    .io_fw_bottom(cells_2d_18_io_fw_bottom),
    .io_fw_right(cells_2d_18_io_fw_right),
    .io_sel(cells_2d_18_io_sel)
  );
  CrossBarCell cells_2d_19 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_19_io_fw_left),
    .io_fw_top(cells_2d_19_io_fw_top),
    .io_fw_bottom(cells_2d_19_io_fw_bottom),
    .io_fw_right(cells_2d_19_io_fw_right),
    .io_sel(cells_2d_19_io_sel)
  );
  CrossBarCell cells_2d_20 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_20_io_fw_left),
    .io_fw_top(cells_2d_20_io_fw_top),
    .io_fw_bottom(cells_2d_20_io_fw_bottom),
    .io_fw_right(cells_2d_20_io_fw_right),
    .io_sel(cells_2d_20_io_sel)
  );
  CrossBarCell cells_2d_21 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_21_io_fw_left),
    .io_fw_top(cells_2d_21_io_fw_top),
    .io_fw_bottom(cells_2d_21_io_fw_bottom),
    .io_fw_right(cells_2d_21_io_fw_right),
    .io_sel(cells_2d_21_io_sel)
  );
  CrossBarCell cells_2d_22 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_22_io_fw_left),
    .io_fw_top(cells_2d_22_io_fw_top),
    .io_fw_bottom(cells_2d_22_io_fw_bottom),
    .io_fw_right(cells_2d_22_io_fw_right),
    .io_sel(cells_2d_22_io_sel)
  );
  CrossBarCell cells_2d_23 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_23_io_fw_left),
    .io_fw_top(cells_2d_23_io_fw_top),
    .io_fw_bottom(cells_2d_23_io_fw_bottom),
    .io_fw_right(cells_2d_23_io_fw_right),
    .io_sel(cells_2d_23_io_sel)
  );
  CrossBarCell cells_2d_24 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_24_io_fw_left),
    .io_fw_top(cells_2d_24_io_fw_top),
    .io_fw_bottom(cells_2d_24_io_fw_bottom),
    .io_fw_right(cells_2d_24_io_fw_right),
    .io_sel(cells_2d_24_io_sel)
  );
  CrossBarCell cells_2d_25 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_25_io_fw_left),
    .io_fw_top(cells_2d_25_io_fw_top),
    .io_fw_bottom(cells_2d_25_io_fw_bottom),
    .io_fw_right(cells_2d_25_io_fw_right),
    .io_sel(cells_2d_25_io_sel)
  );
  CrossBarCell cells_2d_26 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_26_io_fw_left),
    .io_fw_top(cells_2d_26_io_fw_top),
    .io_fw_bottom(cells_2d_26_io_fw_bottom),
    .io_fw_right(cells_2d_26_io_fw_right),
    .io_sel(cells_2d_26_io_sel)
  );
  CrossBarCell cells_2d_27 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_27_io_fw_left),
    .io_fw_top(cells_2d_27_io_fw_top),
    .io_fw_bottom(cells_2d_27_io_fw_bottom),
    .io_fw_right(cells_2d_27_io_fw_right),
    .io_sel(cells_2d_27_io_sel)
  );
  CrossBarCell cells_2d_28 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_28_io_fw_left),
    .io_fw_top(cells_2d_28_io_fw_top),
    .io_fw_bottom(cells_2d_28_io_fw_bottom),
    .io_fw_right(cells_2d_28_io_fw_right),
    .io_sel(cells_2d_28_io_sel)
  );
  CrossBarCell cells_2d_29 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_29_io_fw_left),
    .io_fw_top(cells_2d_29_io_fw_top),
    .io_fw_bottom(cells_2d_29_io_fw_bottom),
    .io_fw_right(cells_2d_29_io_fw_right),
    .io_sel(cells_2d_29_io_sel)
  );
  CrossBarCell cells_2d_30 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_30_io_fw_left),
    .io_fw_top(cells_2d_30_io_fw_top),
    .io_fw_bottom(cells_2d_30_io_fw_bottom),
    .io_fw_right(cells_2d_30_io_fw_right),
    .io_sel(cells_2d_30_io_sel)
  );
  CrossBarCell cells_2d_31 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_31_io_fw_left),
    .io_fw_top(cells_2d_31_io_fw_top),
    .io_fw_bottom(cells_2d_31_io_fw_bottom),
    .io_fw_right(cells_2d_31_io_fw_right),
    .io_sel(cells_2d_31_io_sel)
  );
  CrossBarCell cells_2d_32 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_32_io_fw_left),
    .io_fw_top(cells_2d_32_io_fw_top),
    .io_fw_bottom(cells_2d_32_io_fw_bottom),
    .io_fw_right(cells_2d_32_io_fw_right),
    .io_sel(cells_2d_32_io_sel)
  );
  CrossBarCell cells_2d_33 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_33_io_fw_left),
    .io_fw_top(cells_2d_33_io_fw_top),
    .io_fw_bottom(cells_2d_33_io_fw_bottom),
    .io_fw_right(cells_2d_33_io_fw_right),
    .io_sel(cells_2d_33_io_sel)
  );
  CrossBarCell cells_2d_34 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_34_io_fw_left),
    .io_fw_top(cells_2d_34_io_fw_top),
    .io_fw_bottom(cells_2d_34_io_fw_bottom),
    .io_fw_right(cells_2d_34_io_fw_right),
    .io_sel(cells_2d_34_io_sel)
  );
  CrossBarCell cells_2d_35 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_35_io_fw_left),
    .io_fw_top(cells_2d_35_io_fw_top),
    .io_fw_bottom(cells_2d_35_io_fw_bottom),
    .io_fw_right(cells_2d_35_io_fw_right),
    .io_sel(cells_2d_35_io_sel)
  );
  CrossBarCell cells_2d_36 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_36_io_fw_left),
    .io_fw_top(cells_2d_36_io_fw_top),
    .io_fw_bottom(cells_2d_36_io_fw_bottom),
    .io_fw_right(cells_2d_36_io_fw_right),
    .io_sel(cells_2d_36_io_sel)
  );
  CrossBarCell cells_2d_37 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_37_io_fw_left),
    .io_fw_top(cells_2d_37_io_fw_top),
    .io_fw_bottom(cells_2d_37_io_fw_bottom),
    .io_fw_right(cells_2d_37_io_fw_right),
    .io_sel(cells_2d_37_io_sel)
  );
  CrossBarCell cells_2d_38 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_38_io_fw_left),
    .io_fw_top(cells_2d_38_io_fw_top),
    .io_fw_bottom(cells_2d_38_io_fw_bottom),
    .io_fw_right(cells_2d_38_io_fw_right),
    .io_sel(cells_2d_38_io_sel)
  );
  CrossBarCell cells_2d_39 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_39_io_fw_left),
    .io_fw_top(cells_2d_39_io_fw_top),
    .io_fw_bottom(cells_2d_39_io_fw_bottom),
    .io_fw_right(cells_2d_39_io_fw_right),
    .io_sel(cells_2d_39_io_sel)
  );
  CrossBarCell cells_2d_40 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_40_io_fw_left),
    .io_fw_top(cells_2d_40_io_fw_top),
    .io_fw_bottom(cells_2d_40_io_fw_bottom),
    .io_fw_right(cells_2d_40_io_fw_right),
    .io_sel(cells_2d_40_io_sel)
  );
  CrossBarCell cells_2d_41 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_41_io_fw_left),
    .io_fw_top(cells_2d_41_io_fw_top),
    .io_fw_bottom(cells_2d_41_io_fw_bottom),
    .io_fw_right(cells_2d_41_io_fw_right),
    .io_sel(cells_2d_41_io_sel)
  );
  CrossBarCell cells_2d_42 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_42_io_fw_left),
    .io_fw_top(cells_2d_42_io_fw_top),
    .io_fw_bottom(cells_2d_42_io_fw_bottom),
    .io_fw_right(cells_2d_42_io_fw_right),
    .io_sel(cells_2d_42_io_sel)
  );
  CrossBarCell cells_2d_43 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_43_io_fw_left),
    .io_fw_top(cells_2d_43_io_fw_top),
    .io_fw_bottom(cells_2d_43_io_fw_bottom),
    .io_fw_right(cells_2d_43_io_fw_right),
    .io_sel(cells_2d_43_io_sel)
  );
  CrossBarCell cells_2d_44 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_44_io_fw_left),
    .io_fw_top(cells_2d_44_io_fw_top),
    .io_fw_bottom(cells_2d_44_io_fw_bottom),
    .io_fw_right(cells_2d_44_io_fw_right),
    .io_sel(cells_2d_44_io_sel)
  );
  CrossBarCell cells_2d_45 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_45_io_fw_left),
    .io_fw_top(cells_2d_45_io_fw_top),
    .io_fw_bottom(cells_2d_45_io_fw_bottom),
    .io_fw_right(cells_2d_45_io_fw_right),
    .io_sel(cells_2d_45_io_sel)
  );
  CrossBarCell cells_2d_46 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_46_io_fw_left),
    .io_fw_top(cells_2d_46_io_fw_top),
    .io_fw_bottom(cells_2d_46_io_fw_bottom),
    .io_fw_right(cells_2d_46_io_fw_right),
    .io_sel(cells_2d_46_io_sel)
  );
  CrossBarCell cells_2d_47 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_47_io_fw_left),
    .io_fw_top(cells_2d_47_io_fw_top),
    .io_fw_bottom(cells_2d_47_io_fw_bottom),
    .io_fw_right(cells_2d_47_io_fw_right),
    .io_sel(cells_2d_47_io_sel)
  );
  CrossBarCell cells_2d_48 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_48_io_fw_left),
    .io_fw_top(cells_2d_48_io_fw_top),
    .io_fw_bottom(cells_2d_48_io_fw_bottom),
    .io_fw_right(cells_2d_48_io_fw_right),
    .io_sel(cells_2d_48_io_sel)
  );
  CrossBarCell cells_2d_49 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_49_io_fw_left),
    .io_fw_top(cells_2d_49_io_fw_top),
    .io_fw_bottom(cells_2d_49_io_fw_bottom),
    .io_fw_right(cells_2d_49_io_fw_right),
    .io_sel(cells_2d_49_io_sel)
  );
  CrossBarCell cells_2d_50 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_50_io_fw_left),
    .io_fw_top(cells_2d_50_io_fw_top),
    .io_fw_bottom(cells_2d_50_io_fw_bottom),
    .io_fw_right(cells_2d_50_io_fw_right),
    .io_sel(cells_2d_50_io_sel)
  );
  CrossBarCell cells_2d_51 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_51_io_fw_left),
    .io_fw_top(cells_2d_51_io_fw_top),
    .io_fw_bottom(cells_2d_51_io_fw_bottom),
    .io_fw_right(cells_2d_51_io_fw_right),
    .io_sel(cells_2d_51_io_sel)
  );
  CrossBarCell cells_2d_52 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_52_io_fw_left),
    .io_fw_top(cells_2d_52_io_fw_top),
    .io_fw_bottom(cells_2d_52_io_fw_bottom),
    .io_fw_right(cells_2d_52_io_fw_right),
    .io_sel(cells_2d_52_io_sel)
  );
  CrossBarCell cells_2d_53 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_53_io_fw_left),
    .io_fw_top(cells_2d_53_io_fw_top),
    .io_fw_bottom(cells_2d_53_io_fw_bottom),
    .io_fw_right(cells_2d_53_io_fw_right),
    .io_sel(cells_2d_53_io_sel)
  );
  CrossBarCell cells_2d_54 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_54_io_fw_left),
    .io_fw_top(cells_2d_54_io_fw_top),
    .io_fw_bottom(cells_2d_54_io_fw_bottom),
    .io_fw_right(cells_2d_54_io_fw_right),
    .io_sel(cells_2d_54_io_sel)
  );
  CrossBarCell cells_2d_55 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_55_io_fw_left),
    .io_fw_top(cells_2d_55_io_fw_top),
    .io_fw_bottom(cells_2d_55_io_fw_bottom),
    .io_fw_right(cells_2d_55_io_fw_right),
    .io_sel(cells_2d_55_io_sel)
  );
  CrossBarCell cells_2d_56 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_56_io_fw_left),
    .io_fw_top(cells_2d_56_io_fw_top),
    .io_fw_bottom(cells_2d_56_io_fw_bottom),
    .io_fw_right(cells_2d_56_io_fw_right),
    .io_sel(cells_2d_56_io_sel)
  );
  CrossBarCell cells_2d_57 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_57_io_fw_left),
    .io_fw_top(cells_2d_57_io_fw_top),
    .io_fw_bottom(cells_2d_57_io_fw_bottom),
    .io_fw_right(cells_2d_57_io_fw_right),
    .io_sel(cells_2d_57_io_sel)
  );
  CrossBarCell cells_2d_58 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_58_io_fw_left),
    .io_fw_top(cells_2d_58_io_fw_top),
    .io_fw_bottom(cells_2d_58_io_fw_bottom),
    .io_fw_right(cells_2d_58_io_fw_right),
    .io_sel(cells_2d_58_io_sel)
  );
  CrossBarCell cells_2d_59 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_59_io_fw_left),
    .io_fw_top(cells_2d_59_io_fw_top),
    .io_fw_bottom(cells_2d_59_io_fw_bottom),
    .io_fw_right(cells_2d_59_io_fw_right),
    .io_sel(cells_2d_59_io_sel)
  );
  CrossBarCell cells_2d_60 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_60_io_fw_left),
    .io_fw_top(cells_2d_60_io_fw_top),
    .io_fw_bottom(cells_2d_60_io_fw_bottom),
    .io_fw_right(cells_2d_60_io_fw_right),
    .io_sel(cells_2d_60_io_sel)
  );
  CrossBarCell cells_2d_61 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_61_io_fw_left),
    .io_fw_top(cells_2d_61_io_fw_top),
    .io_fw_bottom(cells_2d_61_io_fw_bottom),
    .io_fw_right(cells_2d_61_io_fw_right),
    .io_sel(cells_2d_61_io_sel)
  );
  CrossBarCell cells_2d_62 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_62_io_fw_left),
    .io_fw_top(cells_2d_62_io_fw_top),
    .io_fw_bottom(cells_2d_62_io_fw_bottom),
    .io_fw_right(cells_2d_62_io_fw_right),
    .io_sel(cells_2d_62_io_sel)
  );
  CrossBarCell cells_2d_63 ( // @[CrossBarSwitchNew.scala 38:53]
    .io_fw_left(cells_2d_63_io_fw_left),
    .io_fw_top(cells_2d_63_io_fw_top),
    .io_fw_bottom(cells_2d_63_io_fw_bottom),
    .io_fw_right(cells_2d_63_io_fw_right),
    .io_sel(cells_2d_63_io_sel)
  );
  assign io_fw_bottom_0 = cells_2d_56_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_1 = cells_2d_57_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_2 = cells_2d_58_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_3 = cells_2d_59_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_4 = cells_2d_60_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_5 = cells_2d_61_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_6 = cells_2d_62_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign io_fw_bottom_7 = cells_2d_63_io_fw_bottom; // @[CrossBarSwitchNew.scala 77:21]
  assign cells_2d_0_io_fw_left = io_fw_left_0; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_0_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_0_io_sel = select_onehot_0[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_1_io_fw_left = cells_2d_0_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_1_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_1_io_sel = select_onehot_1[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_2_io_fw_left = cells_2d_1_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_2_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_2_io_sel = select_onehot_2[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_3_io_fw_left = cells_2d_2_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_3_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_3_io_sel = select_onehot_3[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_4_io_fw_left = cells_2d_3_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_4_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_4_io_sel = select_onehot_4[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_5_io_fw_left = cells_2d_4_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_5_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_5_io_sel = select_onehot_5[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_6_io_fw_left = cells_2d_5_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_6_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_6_io_sel = select_onehot_6[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_7_io_fw_left = cells_2d_6_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_7_io_fw_top = 64'h0; // @[CrossBarSwitchNew.scala 56:28]
  assign cells_2d_7_io_sel = select_onehot_7[0]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_8_io_fw_left = io_fw_left_1; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_8_io_fw_top = cells_2d_0_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_8_io_sel = select_onehot_0[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_9_io_fw_left = cells_2d_8_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_9_io_fw_top = cells_2d_1_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_9_io_sel = select_onehot_1[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_10_io_fw_left = cells_2d_9_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_10_io_fw_top = cells_2d_2_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_10_io_sel = select_onehot_2[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_11_io_fw_left = cells_2d_10_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_11_io_fw_top = cells_2d_3_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_11_io_sel = select_onehot_3[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_12_io_fw_left = cells_2d_11_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_12_io_fw_top = cells_2d_4_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_12_io_sel = select_onehot_4[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_13_io_fw_left = cells_2d_12_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_13_io_fw_top = cells_2d_5_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_13_io_sel = select_onehot_5[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_14_io_fw_left = cells_2d_13_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_14_io_fw_top = cells_2d_6_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_14_io_sel = select_onehot_6[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_15_io_fw_left = cells_2d_14_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_15_io_fw_top = cells_2d_7_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_15_io_sel = select_onehot_7[1]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_16_io_fw_left = io_fw_left_2; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_16_io_fw_top = cells_2d_8_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_16_io_sel = select_onehot_0[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_17_io_fw_left = cells_2d_16_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_17_io_fw_top = cells_2d_9_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_17_io_sel = select_onehot_1[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_18_io_fw_left = cells_2d_17_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_18_io_fw_top = cells_2d_10_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_18_io_sel = select_onehot_2[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_19_io_fw_left = cells_2d_18_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_19_io_fw_top = cells_2d_11_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_19_io_sel = select_onehot_3[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_20_io_fw_left = cells_2d_19_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_20_io_fw_top = cells_2d_12_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_20_io_sel = select_onehot_4[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_21_io_fw_left = cells_2d_20_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_21_io_fw_top = cells_2d_13_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_21_io_sel = select_onehot_5[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_22_io_fw_left = cells_2d_21_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_22_io_fw_top = cells_2d_14_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_22_io_sel = select_onehot_6[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_23_io_fw_left = cells_2d_22_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_23_io_fw_top = cells_2d_15_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_23_io_sel = select_onehot_7[2]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_24_io_fw_left = io_fw_left_3; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_24_io_fw_top = cells_2d_16_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_24_io_sel = select_onehot_0[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_25_io_fw_left = cells_2d_24_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_25_io_fw_top = cells_2d_17_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_25_io_sel = select_onehot_1[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_26_io_fw_left = cells_2d_25_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_26_io_fw_top = cells_2d_18_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_26_io_sel = select_onehot_2[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_27_io_fw_left = cells_2d_26_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_27_io_fw_top = cells_2d_19_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_27_io_sel = select_onehot_3[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_28_io_fw_left = cells_2d_27_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_28_io_fw_top = cells_2d_20_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_28_io_sel = select_onehot_4[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_29_io_fw_left = cells_2d_28_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_29_io_fw_top = cells_2d_21_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_29_io_sel = select_onehot_5[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_30_io_fw_left = cells_2d_29_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_30_io_fw_top = cells_2d_22_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_30_io_sel = select_onehot_6[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_31_io_fw_left = cells_2d_30_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_31_io_fw_top = cells_2d_23_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_31_io_sel = select_onehot_7[3]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_32_io_fw_left = io_fw_left_4; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_32_io_fw_top = cells_2d_24_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_32_io_sel = select_onehot_0[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_33_io_fw_left = cells_2d_32_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_33_io_fw_top = cells_2d_25_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_33_io_sel = select_onehot_1[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_34_io_fw_left = cells_2d_33_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_34_io_fw_top = cells_2d_26_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_34_io_sel = select_onehot_2[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_35_io_fw_left = cells_2d_34_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_35_io_fw_top = cells_2d_27_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_35_io_sel = select_onehot_3[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_36_io_fw_left = cells_2d_35_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_36_io_fw_top = cells_2d_28_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_36_io_sel = select_onehot_4[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_37_io_fw_left = cells_2d_36_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_37_io_fw_top = cells_2d_29_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_37_io_sel = select_onehot_5[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_38_io_fw_left = cells_2d_37_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_38_io_fw_top = cells_2d_30_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_38_io_sel = select_onehot_6[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_39_io_fw_left = cells_2d_38_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_39_io_fw_top = cells_2d_31_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_39_io_sel = select_onehot_7[4]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_40_io_fw_left = io_fw_left_5; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_40_io_fw_top = cells_2d_32_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_40_io_sel = select_onehot_0[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_41_io_fw_left = cells_2d_40_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_41_io_fw_top = cells_2d_33_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_41_io_sel = select_onehot_1[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_42_io_fw_left = cells_2d_41_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_42_io_fw_top = cells_2d_34_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_42_io_sel = select_onehot_2[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_43_io_fw_left = cells_2d_42_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_43_io_fw_top = cells_2d_35_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_43_io_sel = select_onehot_3[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_44_io_fw_left = cells_2d_43_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_44_io_fw_top = cells_2d_36_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_44_io_sel = select_onehot_4[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_45_io_fw_left = cells_2d_44_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_45_io_fw_top = cells_2d_37_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_45_io_sel = select_onehot_5[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_46_io_fw_left = cells_2d_45_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_46_io_fw_top = cells_2d_38_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_46_io_sel = select_onehot_6[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_47_io_fw_left = cells_2d_46_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_47_io_fw_top = cells_2d_39_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_47_io_sel = select_onehot_7[5]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_48_io_fw_left = io_fw_left_6; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_48_io_fw_top = cells_2d_40_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_48_io_sel = select_onehot_0[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_49_io_fw_left = cells_2d_48_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_49_io_fw_top = cells_2d_41_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_49_io_sel = select_onehot_1[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_50_io_fw_left = cells_2d_49_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_50_io_fw_top = cells_2d_42_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_50_io_sel = select_onehot_2[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_51_io_fw_left = cells_2d_50_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_51_io_fw_top = cells_2d_43_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_51_io_sel = select_onehot_3[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_52_io_fw_left = cells_2d_51_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_52_io_fw_top = cells_2d_44_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_52_io_sel = select_onehot_4[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_53_io_fw_left = cells_2d_52_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_53_io_fw_top = cells_2d_45_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_53_io_sel = select_onehot_5[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_54_io_fw_left = cells_2d_53_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_54_io_fw_top = cells_2d_46_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_54_io_sel = select_onehot_6[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_55_io_fw_left = cells_2d_54_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_55_io_fw_top = cells_2d_47_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_55_io_sel = select_onehot_7[6]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_56_io_fw_left = io_fw_left_7; // @[CrossBarSwitchNew.scala 63:29]
  assign cells_2d_56_io_fw_top = cells_2d_48_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_56_io_sel = select_onehot_0[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_57_io_fw_left = cells_2d_56_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_57_io_fw_top = cells_2d_49_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_57_io_sel = select_onehot_1[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_58_io_fw_left = cells_2d_57_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_58_io_fw_top = cells_2d_50_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_58_io_sel = select_onehot_2[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_59_io_fw_left = cells_2d_58_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_59_io_fw_top = cells_2d_51_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_59_io_sel = select_onehot_3[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_60_io_fw_left = cells_2d_59_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_60_io_fw_top = cells_2d_52_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_60_io_sel = select_onehot_4[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_61_io_fw_left = cells_2d_60_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_61_io_fw_top = cells_2d_53_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_61_io_sel = select_onehot_5[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_62_io_fw_left = cells_2d_61_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_62_io_fw_top = cells_2d_54_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_62_io_sel = select_onehot_6[7]; // @[CrossBarSwitchNew.scala 70:44]
  assign cells_2d_63_io_fw_left = cells_2d_62_io_fw_right; // @[CrossBarSwitchNew.scala 66:29]
  assign cells_2d_63_io_fw_top = cells_2d_55_io_fw_bottom; // @[CrossBarSwitchNew.scala 59:28]
  assign cells_2d_63_io_sel = select_onehot_7[7]; // @[CrossBarSwitchNew.scala 70:44]
endmodule
module RegMux(
  input         clock,
  input  [63:0] io_in,
  output [63:0] io_out,
  input         io_sel
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] reg_; // @[RegMux.scala 11:16]
  wire [63:0] _GEN_0 = io_sel ? reg_ : io_in; // @[RegMux.scala 15:32 RegMux.scala 16:12 RegMux.scala 18:12]
  assign io_out = ~io_sel ? io_in : _GEN_0; // @[RegMux.scala 13:27 RegMux.scala 14:12]
  always @(posedge clock) begin
    reg_ <= io_in; // @[RegMux.scala 12:7]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  reg_ = _RAND_0[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Tile(
  input         clock,
  input         reset,
  input  [31:0] io_controlSignal_wr,
  input         io_controlSignal_wr_en,
  input         io_run,
  input  [63:0] io_north_in_a,
  input  [63:0] io_north_in_b,
  output [63:0] io_north_out_a,
  output [63:0] io_north_out_b,
  input  [63:0] io_east_in_a,
  input  [63:0] io_east_in_b,
  output [63:0] io_east_out_a,
  output [63:0] io_east_out_b,
  input  [63:0] io_west_in_a,
  input  [63:0] io_west_in_b,
  output [63:0] io_west_out_a,
  output [63:0] io_west_out_b,
  input  [63:0] io_south_in_a,
  input  [63:0] io_south_in_b,
  output [63:0] io_south_out_a,
  output [63:0] io_south_out_b
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mem [0:1023]; // @[Tile.scala 54:16]
  wire [63:0] mem_ctrl_MPORT_data; // @[Tile.scala 54:16]
  wire [9:0] mem_ctrl_MPORT_addr; // @[Tile.scala 54:16]
  wire [63:0] mem_MPORT_data; // @[Tile.scala 54:16]
  wire [9:0] mem_MPORT_addr; // @[Tile.scala 54:16]
  wire  mem_MPORT_mask; // @[Tile.scala 54:16]
  wire  mem_MPORT_en; // @[Tile.scala 54:16]
  wire [63:0] crossBar_io_fw_left_0; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_left_1; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_left_2; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_left_3; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_left_4; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_left_5; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_left_6; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_left_7; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_0; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_1; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_2; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_3; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_4; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_5; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_6; // @[Tile.scala 70:24]
  wire [63:0] crossBar_io_fw_bottom_7; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_0; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_1; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_2; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_3; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_4; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_5; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_6; // @[Tile.scala 70:24]
  wire [2:0] crossBar_io_select_7; // @[Tile.scala 70:24]
  wire  RegMux_clock; // @[Tile.scala 90:59]
  wire [63:0] RegMux_io_in; // @[Tile.scala 90:59]
  wire [63:0] RegMux_io_out; // @[Tile.scala 90:59]
  wire  RegMux_io_sel; // @[Tile.scala 90:59]
  wire  RegMux_1_clock; // @[Tile.scala 90:59]
  wire [63:0] RegMux_1_io_in; // @[Tile.scala 90:59]
  wire [63:0] RegMux_1_io_out; // @[Tile.scala 90:59]
  wire  RegMux_1_io_sel; // @[Tile.scala 90:59]
  wire  RegMux_2_clock; // @[Tile.scala 102:58]
  wire [63:0] RegMux_2_io_in; // @[Tile.scala 102:58]
  wire [63:0] RegMux_2_io_out; // @[Tile.scala 102:58]
  wire  RegMux_2_io_sel; // @[Tile.scala 102:58]
  wire  RegMux_3_clock; // @[Tile.scala 102:58]
  wire [63:0] RegMux_3_io_in; // @[Tile.scala 102:58]
  wire [63:0] RegMux_3_io_out; // @[Tile.scala 102:58]
  wire  RegMux_3_io_sel; // @[Tile.scala 102:58]
  wire  RegMux_4_clock; // @[Tile.scala 114:58]
  wire [63:0] RegMux_4_io_in; // @[Tile.scala 114:58]
  wire [63:0] RegMux_4_io_out; // @[Tile.scala 114:58]
  wire  RegMux_4_io_sel; // @[Tile.scala 114:58]
  wire  RegMux_5_clock; // @[Tile.scala 114:58]
  wire [63:0] RegMux_5_io_in; // @[Tile.scala 114:58]
  wire [63:0] RegMux_5_io_out; // @[Tile.scala 114:58]
  wire  RegMux_5_io_sel; // @[Tile.scala 114:58]
  wire  RegMux_6_clock; // @[Tile.scala 126:59]
  wire [63:0] RegMux_6_io_in; // @[Tile.scala 126:59]
  wire [63:0] RegMux_6_io_out; // @[Tile.scala 126:59]
  wire  RegMux_6_io_sel; // @[Tile.scala 126:59]
  wire  RegMux_7_clock; // @[Tile.scala 126:59]
  wire [63:0] RegMux_7_io_in; // @[Tile.scala 126:59]
  wire [63:0] RegMux_7_io_out; // @[Tile.scala 126:59]
  wire  RegMux_7_io_sel; // @[Tile.scala 126:59]
  reg [9:0] rdAddrBase; // @[Tile.scala 55:27]
  reg [9:0] wrAddrBase; // @[Tile.scala 56:27]
  reg [63:0] ctrl; // @[Tile.scala 57:21]
  wire [9:0] _wrAddrBase_T_1 = wrAddrBase + 10'h1; // @[Tile.scala 61:30]
  wire [9:0] _rdAddrBase_T_1 = rdAddrBase + 10'h1; // @[Tile.scala 66:30]
  wire [7:0] RegMuxSel = ctrl[36:29]; // @[Tile.scala 73:23]
  wire [23:0] CrossBarSel = ctrl[28:5]; // @[Tile.scala 74:25]
  CrossBarSwitchNew crossBar ( // @[Tile.scala 70:24]
    .io_fw_left_0(crossBar_io_fw_left_0),
    .io_fw_left_1(crossBar_io_fw_left_1),
    .io_fw_left_2(crossBar_io_fw_left_2),
    .io_fw_left_3(crossBar_io_fw_left_3),
    .io_fw_left_4(crossBar_io_fw_left_4),
    .io_fw_left_5(crossBar_io_fw_left_5),
    .io_fw_left_6(crossBar_io_fw_left_6),
    .io_fw_left_7(crossBar_io_fw_left_7),
    .io_fw_bottom_0(crossBar_io_fw_bottom_0),
    .io_fw_bottom_1(crossBar_io_fw_bottom_1),
    .io_fw_bottom_2(crossBar_io_fw_bottom_2),
    .io_fw_bottom_3(crossBar_io_fw_bottom_3),
    .io_fw_bottom_4(crossBar_io_fw_bottom_4),
    .io_fw_bottom_5(crossBar_io_fw_bottom_5),
    .io_fw_bottom_6(crossBar_io_fw_bottom_6),
    .io_fw_bottom_7(crossBar_io_fw_bottom_7),
    .io_select_0(crossBar_io_select_0),
    .io_select_1(crossBar_io_select_1),
    .io_select_2(crossBar_io_select_2),
    .io_select_3(crossBar_io_select_3),
    .io_select_4(crossBar_io_select_4),
    .io_select_5(crossBar_io_select_5),
    .io_select_6(crossBar_io_select_6),
    .io_select_7(crossBar_io_select_7)
  );
  RegMux RegMux ( // @[Tile.scala 90:59]
    .clock(RegMux_clock),
    .io_in(RegMux_io_in),
    .io_out(RegMux_io_out),
    .io_sel(RegMux_io_sel)
  );
  RegMux RegMux_1 ( // @[Tile.scala 90:59]
    .clock(RegMux_1_clock),
    .io_in(RegMux_1_io_in),
    .io_out(RegMux_1_io_out),
    .io_sel(RegMux_1_io_sel)
  );
  RegMux RegMux_2 ( // @[Tile.scala 102:58]
    .clock(RegMux_2_clock),
    .io_in(RegMux_2_io_in),
    .io_out(RegMux_2_io_out),
    .io_sel(RegMux_2_io_sel)
  );
  RegMux RegMux_3 ( // @[Tile.scala 102:58]
    .clock(RegMux_3_clock),
    .io_in(RegMux_3_io_in),
    .io_out(RegMux_3_io_out),
    .io_sel(RegMux_3_io_sel)
  );
  RegMux RegMux_4 ( // @[Tile.scala 114:58]
    .clock(RegMux_4_clock),
    .io_in(RegMux_4_io_in),
    .io_out(RegMux_4_io_out),
    .io_sel(RegMux_4_io_sel)
  );
  RegMux RegMux_5 ( // @[Tile.scala 114:58]
    .clock(RegMux_5_clock),
    .io_in(RegMux_5_io_in),
    .io_out(RegMux_5_io_out),
    .io_sel(RegMux_5_io_sel)
  );
  RegMux RegMux_6 ( // @[Tile.scala 126:59]
    .clock(RegMux_6_clock),
    .io_in(RegMux_6_io_in),
    .io_out(RegMux_6_io_out),
    .io_sel(RegMux_6_io_sel)
  );
  RegMux RegMux_7 ( // @[Tile.scala 126:59]
    .clock(RegMux_7_clock),
    .io_in(RegMux_7_io_in),
    .io_out(RegMux_7_io_out),
    .io_sel(RegMux_7_io_sel)
  );
  assign mem_ctrl_MPORT_addr = rdAddrBase;
  assign mem_ctrl_MPORT_data = mem[mem_ctrl_MPORT_addr]; // @[Tile.scala 54:16]
  assign mem_MPORT_data = {{32'd0}, io_controlSignal_wr};
  assign mem_MPORT_addr = wrAddrBase;
  assign mem_MPORT_mask = 1'h1;
  assign mem_MPORT_en = io_controlSignal_wr_en;
  assign io_north_out_a = crossBar_io_fw_bottom_0; // @[Tile.scala 136:18]
  assign io_north_out_b = crossBar_io_fw_bottom_1; // @[Tile.scala 137:18]
  assign io_east_out_a = crossBar_io_fw_bottom_2; // @[Tile.scala 138:17]
  assign io_east_out_b = crossBar_io_fw_bottom_3; // @[Tile.scala 139:17]
  assign io_west_out_a = crossBar_io_fw_bottom_4; // @[Tile.scala 140:17]
  assign io_west_out_b = crossBar_io_fw_bottom_5; // @[Tile.scala 141:17]
  assign io_south_out_a = crossBar_io_fw_bottom_6; // @[Tile.scala 142:18]
  assign io_south_out_b = crossBar_io_fw_bottom_7; // @[Tile.scala 143:18]
  assign crossBar_io_fw_left_0 = RegMux_io_out; // @[Tile.scala 93:28]
  assign crossBar_io_fw_left_1 = RegMux_1_io_out; // @[Tile.scala 97:28]
  assign crossBar_io_fw_left_2 = RegMux_2_io_out; // @[Tile.scala 105:28]
  assign crossBar_io_fw_left_3 = RegMux_3_io_out; // @[Tile.scala 109:28]
  assign crossBar_io_fw_left_4 = RegMux_4_io_out; // @[Tile.scala 117:28]
  assign crossBar_io_fw_left_5 = RegMux_5_io_out; // @[Tile.scala 121:28]
  assign crossBar_io_fw_left_6 = RegMux_6_io_out; // @[Tile.scala 129:28]
  assign crossBar_io_fw_left_7 = RegMux_7_io_out; // @[Tile.scala 133:28]
  assign crossBar_io_select_0 = CrossBarSel[2:0]; // @[Tile.scala 81:37]
  assign crossBar_io_select_1 = CrossBarSel[5:3]; // @[Tile.scala 81:37]
  assign crossBar_io_select_2 = CrossBarSel[8:6]; // @[Tile.scala 81:37]
  assign crossBar_io_select_3 = CrossBarSel[11:9]; // @[Tile.scala 81:37]
  assign crossBar_io_select_4 = CrossBarSel[14:12]; // @[Tile.scala 81:37]
  assign crossBar_io_select_5 = CrossBarSel[17:15]; // @[Tile.scala 81:37]
  assign crossBar_io_select_6 = CrossBarSel[20:18]; // @[Tile.scala 81:37]
  assign crossBar_io_select_7 = CrossBarSel[23:21]; // @[Tile.scala 81:37]
  assign RegMux_clock = clock;
  assign RegMux_io_in = io_north_in_a; // @[Tile.scala 91:26]
  assign RegMux_io_sel = RegMuxSel[0]; // @[Tile.scala 92:45]
  assign RegMux_1_clock = clock;
  assign RegMux_1_io_in = io_north_in_b; // @[Tile.scala 95:26]
  assign RegMux_1_io_sel = RegMuxSel[1]; // @[Tile.scala 96:45]
  assign RegMux_2_clock = clock;
  assign RegMux_2_io_in = io_east_in_a; // @[Tile.scala 103:25]
  assign RegMux_2_io_sel = RegMuxSel[2]; // @[Tile.scala 104:44]
  assign RegMux_3_clock = clock;
  assign RegMux_3_io_in = io_east_in_b; // @[Tile.scala 107:25]
  assign RegMux_3_io_sel = RegMuxSel[3]; // @[Tile.scala 108:44]
  assign RegMux_4_clock = clock;
  assign RegMux_4_io_in = io_west_in_a; // @[Tile.scala 115:25]
  assign RegMux_4_io_sel = RegMuxSel[4]; // @[Tile.scala 116:44]
  assign RegMux_5_clock = clock;
  assign RegMux_5_io_in = io_west_in_b; // @[Tile.scala 119:25]
  assign RegMux_5_io_sel = RegMuxSel[5]; // @[Tile.scala 120:44]
  assign RegMux_6_clock = clock;
  assign RegMux_6_io_in = io_south_in_a; // @[Tile.scala 127:26]
  assign RegMux_6_io_sel = RegMuxSel[6]; // @[Tile.scala 128:45]
  assign RegMux_7_clock = clock;
  assign RegMux_7_io_in = io_south_in_b; // @[Tile.scala 131:26]
  assign RegMux_7_io_sel = RegMuxSel[7]; // @[Tile.scala 132:45]
  always @(posedge clock) begin
    if(mem_MPORT_en & mem_MPORT_mask) begin
      mem[mem_MPORT_addr] <= mem_MPORT_data; // @[Tile.scala 54:16]
    end
    if (reset) begin // @[Tile.scala 55:27]
      rdAddrBase <= 10'h0; // @[Tile.scala 55:27]
    end else if (io_run) begin // @[Tile.scala 64:16]
      rdAddrBase <= _rdAddrBase_T_1; // @[Tile.scala 66:16]
    end
    if (reset) begin // @[Tile.scala 56:27]
      wrAddrBase <= 10'h0; // @[Tile.scala 56:27]
    end else if (io_controlSignal_wr_en) begin // @[Tile.scala 59:32]
      wrAddrBase <= _wrAddrBase_T_1; // @[Tile.scala 61:16]
    end
    if (reset) begin // @[Tile.scala 57:21]
      ctrl <= 64'h0; // @[Tile.scala 57:21]
    end else if (io_run) begin // @[Tile.scala 64:16]
      ctrl <= mem_ctrl_MPORT_data; // @[Tile.scala 65:10]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    mem[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rdAddrBase = _RAND_1[9:0];
  _RAND_2 = {1{`RANDOM}};
  wrAddrBase = _RAND_2[9:0];
  _RAND_3 = {2{`RANDOM}};
  ctrl = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
