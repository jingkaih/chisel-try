module CrossBarCell(
  input  [63:0] io_fw_left,
  input  [63:0] io_fw_top,
  output [63:0] io_fw_bottom,
  output [63:0] io_fw_right,
  input         io_sel
);
  assign io_fw_bottom = io_sel ? io_fw_left : io_fw_top; // @[CrossBarSwitch.scala 15:17 CrossBarSwitch.scala 16:18 CrossBarSwitch.scala 18:18]
  assign io_fw_right = io_fw_left; // @[CrossBarSwitch.scala 14:15]
endmodule
module CrossBarSwitch(
  input         clock,
  input         reset,
  input  [63:0] io_fw_left_0,
  input  [63:0] io_fw_left_1,
  input  [63:0] io_fw_left_2,
  input  [63:0] io_fw_left_3,
  input  [63:0] io_fw_left_4,
  input  [63:0] io_fw_left_5,
  input  [63:0] io_fw_left_6,
  input  [63:0] io_fw_left_7,
  output [63:0] io_fw_bottom_0,
  output [63:0] io_fw_bottom_1,
  output [63:0] io_fw_bottom_2,
  output [63:0] io_fw_bottom_3,
  output [63:0] io_fw_bottom_4,
  output [63:0] io_fw_bottom_5,
  output [63:0] io_fw_bottom_6,
  output [63:0] io_fw_bottom_7,
  input  [2:0]  io_select_0,
  input  [2:0]  io_select_1,
  input  [2:0]  io_select_2,
  input  [2:0]  io_select_3,
  input  [2:0]  io_select_4,
  input  [2:0]  io_select_5,
  input  [2:0]  io_select_6,
  input  [2:0]  io_select_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [63:0] cells_2d_0_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_0_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_0_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_0_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_0_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_1_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_1_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_1_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_1_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_1_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_2_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_2_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_2_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_2_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_2_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_3_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_3_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_3_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_3_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_3_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_4_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_4_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_4_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_4_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_4_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_5_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_5_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_5_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_5_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_5_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_6_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_6_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_6_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_6_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_6_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_7_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_7_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_7_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_7_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_7_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_8_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_8_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_8_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_8_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_8_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_9_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_9_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_9_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_9_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_9_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_10_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_10_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_10_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_10_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_10_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_11_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_11_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_11_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_11_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_11_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_12_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_12_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_12_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_12_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_12_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_13_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_13_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_13_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_13_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_13_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_14_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_14_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_14_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_14_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_14_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_15_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_15_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_15_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_15_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_15_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_16_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_16_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_16_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_16_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_16_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_17_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_17_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_17_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_17_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_17_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_18_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_18_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_18_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_18_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_18_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_19_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_19_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_19_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_19_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_19_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_20_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_20_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_20_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_20_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_20_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_21_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_21_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_21_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_21_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_21_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_22_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_22_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_22_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_22_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_22_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_23_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_23_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_23_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_23_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_23_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_24_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_24_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_24_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_24_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_24_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_25_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_25_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_25_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_25_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_25_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_26_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_26_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_26_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_26_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_26_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_27_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_27_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_27_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_27_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_27_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_28_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_28_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_28_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_28_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_28_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_29_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_29_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_29_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_29_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_29_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_30_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_30_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_30_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_30_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_30_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_31_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_31_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_31_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_31_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_31_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_32_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_32_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_32_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_32_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_32_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_33_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_33_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_33_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_33_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_33_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_34_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_34_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_34_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_34_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_34_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_35_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_35_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_35_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_35_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_35_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_36_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_36_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_36_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_36_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_36_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_37_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_37_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_37_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_37_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_37_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_38_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_38_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_38_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_38_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_38_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_39_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_39_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_39_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_39_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_39_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_40_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_40_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_40_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_40_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_40_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_41_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_41_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_41_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_41_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_41_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_42_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_42_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_42_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_42_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_42_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_43_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_43_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_43_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_43_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_43_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_44_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_44_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_44_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_44_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_44_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_45_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_45_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_45_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_45_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_45_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_46_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_46_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_46_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_46_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_46_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_47_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_47_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_47_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_47_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_47_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_48_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_48_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_48_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_48_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_48_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_49_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_49_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_49_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_49_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_49_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_50_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_50_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_50_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_50_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_50_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_51_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_51_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_51_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_51_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_51_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_52_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_52_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_52_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_52_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_52_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_53_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_53_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_53_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_53_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_53_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_54_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_54_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_54_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_54_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_54_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_55_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_55_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_55_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_55_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_55_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_56_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_56_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_56_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_56_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_56_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_57_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_57_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_57_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_57_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_57_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_58_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_58_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_58_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_58_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_58_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_59_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_59_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_59_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_59_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_59_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_60_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_60_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_60_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_60_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_60_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_61_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_61_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_61_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_61_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_61_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_62_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_62_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_62_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_62_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_62_io_sel; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_63_io_fw_left; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_63_io_fw_top; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_63_io_fw_bottom; // @[CrossBarSwitch.scala 37:53]
  wire [63:0] cells_2d_63_io_fw_right; // @[CrossBarSwitch.scala 37:53]
  wire  cells_2d_63_io_sel; // @[CrossBarSwitch.scala 37:53]
  reg [63:0] fw_left_reg_0; // @[CrossBarSwitch.scala 33:28]
  reg [63:0] fw_left_reg_1; // @[CrossBarSwitch.scala 33:28]
  reg [63:0] fw_left_reg_2; // @[CrossBarSwitch.scala 33:28]
  reg [63:0] fw_left_reg_3; // @[CrossBarSwitch.scala 33:28]
  reg [63:0] fw_left_reg_4; // @[CrossBarSwitch.scala 33:28]
  reg [63:0] fw_left_reg_5; // @[CrossBarSwitch.scala 33:28]
  reg [63:0] fw_left_reg_6; // @[CrossBarSwitch.scala 33:28]
  reg [63:0] fw_left_reg_7; // @[CrossBarSwitch.scala 33:28]
  wire [7:0] select_onehot_0 = 8'h1 << io_select_0; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_1 = 8'h1 << io_select_1; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_2 = 8'h1 << io_select_2; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_3 = 8'h1 << io_select_3; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_4 = 8'h1 << io_select_4; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_5 = 8'h1 << io_select_5; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_6 = 8'h1 << io_select_6; // @[OneHot.scala 65:12]
  wire [7:0] select_onehot_7 = 8'h1 << io_select_7; // @[OneHot.scala 65:12]
  CrossBarCell cells_2d_0 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_0_io_fw_left),
    .io_fw_top(cells_2d_0_io_fw_top),
    .io_fw_bottom(cells_2d_0_io_fw_bottom),
    .io_fw_right(cells_2d_0_io_fw_right),
    .io_sel(cells_2d_0_io_sel)
  );
  CrossBarCell cells_2d_1 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_1_io_fw_left),
    .io_fw_top(cells_2d_1_io_fw_top),
    .io_fw_bottom(cells_2d_1_io_fw_bottom),
    .io_fw_right(cells_2d_1_io_fw_right),
    .io_sel(cells_2d_1_io_sel)
  );
  CrossBarCell cells_2d_2 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_2_io_fw_left),
    .io_fw_top(cells_2d_2_io_fw_top),
    .io_fw_bottom(cells_2d_2_io_fw_bottom),
    .io_fw_right(cells_2d_2_io_fw_right),
    .io_sel(cells_2d_2_io_sel)
  );
  CrossBarCell cells_2d_3 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_3_io_fw_left),
    .io_fw_top(cells_2d_3_io_fw_top),
    .io_fw_bottom(cells_2d_3_io_fw_bottom),
    .io_fw_right(cells_2d_3_io_fw_right),
    .io_sel(cells_2d_3_io_sel)
  );
  CrossBarCell cells_2d_4 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_4_io_fw_left),
    .io_fw_top(cells_2d_4_io_fw_top),
    .io_fw_bottom(cells_2d_4_io_fw_bottom),
    .io_fw_right(cells_2d_4_io_fw_right),
    .io_sel(cells_2d_4_io_sel)
  );
  CrossBarCell cells_2d_5 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_5_io_fw_left),
    .io_fw_top(cells_2d_5_io_fw_top),
    .io_fw_bottom(cells_2d_5_io_fw_bottom),
    .io_fw_right(cells_2d_5_io_fw_right),
    .io_sel(cells_2d_5_io_sel)
  );
  CrossBarCell cells_2d_6 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_6_io_fw_left),
    .io_fw_top(cells_2d_6_io_fw_top),
    .io_fw_bottom(cells_2d_6_io_fw_bottom),
    .io_fw_right(cells_2d_6_io_fw_right),
    .io_sel(cells_2d_6_io_sel)
  );
  CrossBarCell cells_2d_7 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_7_io_fw_left),
    .io_fw_top(cells_2d_7_io_fw_top),
    .io_fw_bottom(cells_2d_7_io_fw_bottom),
    .io_fw_right(cells_2d_7_io_fw_right),
    .io_sel(cells_2d_7_io_sel)
  );
  CrossBarCell cells_2d_8 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_8_io_fw_left),
    .io_fw_top(cells_2d_8_io_fw_top),
    .io_fw_bottom(cells_2d_8_io_fw_bottom),
    .io_fw_right(cells_2d_8_io_fw_right),
    .io_sel(cells_2d_8_io_sel)
  );
  CrossBarCell cells_2d_9 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_9_io_fw_left),
    .io_fw_top(cells_2d_9_io_fw_top),
    .io_fw_bottom(cells_2d_9_io_fw_bottom),
    .io_fw_right(cells_2d_9_io_fw_right),
    .io_sel(cells_2d_9_io_sel)
  );
  CrossBarCell cells_2d_10 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_10_io_fw_left),
    .io_fw_top(cells_2d_10_io_fw_top),
    .io_fw_bottom(cells_2d_10_io_fw_bottom),
    .io_fw_right(cells_2d_10_io_fw_right),
    .io_sel(cells_2d_10_io_sel)
  );
  CrossBarCell cells_2d_11 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_11_io_fw_left),
    .io_fw_top(cells_2d_11_io_fw_top),
    .io_fw_bottom(cells_2d_11_io_fw_bottom),
    .io_fw_right(cells_2d_11_io_fw_right),
    .io_sel(cells_2d_11_io_sel)
  );
  CrossBarCell cells_2d_12 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_12_io_fw_left),
    .io_fw_top(cells_2d_12_io_fw_top),
    .io_fw_bottom(cells_2d_12_io_fw_bottom),
    .io_fw_right(cells_2d_12_io_fw_right),
    .io_sel(cells_2d_12_io_sel)
  );
  CrossBarCell cells_2d_13 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_13_io_fw_left),
    .io_fw_top(cells_2d_13_io_fw_top),
    .io_fw_bottom(cells_2d_13_io_fw_bottom),
    .io_fw_right(cells_2d_13_io_fw_right),
    .io_sel(cells_2d_13_io_sel)
  );
  CrossBarCell cells_2d_14 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_14_io_fw_left),
    .io_fw_top(cells_2d_14_io_fw_top),
    .io_fw_bottom(cells_2d_14_io_fw_bottom),
    .io_fw_right(cells_2d_14_io_fw_right),
    .io_sel(cells_2d_14_io_sel)
  );
  CrossBarCell cells_2d_15 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_15_io_fw_left),
    .io_fw_top(cells_2d_15_io_fw_top),
    .io_fw_bottom(cells_2d_15_io_fw_bottom),
    .io_fw_right(cells_2d_15_io_fw_right),
    .io_sel(cells_2d_15_io_sel)
  );
  CrossBarCell cells_2d_16 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_16_io_fw_left),
    .io_fw_top(cells_2d_16_io_fw_top),
    .io_fw_bottom(cells_2d_16_io_fw_bottom),
    .io_fw_right(cells_2d_16_io_fw_right),
    .io_sel(cells_2d_16_io_sel)
  );
  CrossBarCell cells_2d_17 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_17_io_fw_left),
    .io_fw_top(cells_2d_17_io_fw_top),
    .io_fw_bottom(cells_2d_17_io_fw_bottom),
    .io_fw_right(cells_2d_17_io_fw_right),
    .io_sel(cells_2d_17_io_sel)
  );
  CrossBarCell cells_2d_18 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_18_io_fw_left),
    .io_fw_top(cells_2d_18_io_fw_top),
    .io_fw_bottom(cells_2d_18_io_fw_bottom),
    .io_fw_right(cells_2d_18_io_fw_right),
    .io_sel(cells_2d_18_io_sel)
  );
  CrossBarCell cells_2d_19 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_19_io_fw_left),
    .io_fw_top(cells_2d_19_io_fw_top),
    .io_fw_bottom(cells_2d_19_io_fw_bottom),
    .io_fw_right(cells_2d_19_io_fw_right),
    .io_sel(cells_2d_19_io_sel)
  );
  CrossBarCell cells_2d_20 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_20_io_fw_left),
    .io_fw_top(cells_2d_20_io_fw_top),
    .io_fw_bottom(cells_2d_20_io_fw_bottom),
    .io_fw_right(cells_2d_20_io_fw_right),
    .io_sel(cells_2d_20_io_sel)
  );
  CrossBarCell cells_2d_21 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_21_io_fw_left),
    .io_fw_top(cells_2d_21_io_fw_top),
    .io_fw_bottom(cells_2d_21_io_fw_bottom),
    .io_fw_right(cells_2d_21_io_fw_right),
    .io_sel(cells_2d_21_io_sel)
  );
  CrossBarCell cells_2d_22 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_22_io_fw_left),
    .io_fw_top(cells_2d_22_io_fw_top),
    .io_fw_bottom(cells_2d_22_io_fw_bottom),
    .io_fw_right(cells_2d_22_io_fw_right),
    .io_sel(cells_2d_22_io_sel)
  );
  CrossBarCell cells_2d_23 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_23_io_fw_left),
    .io_fw_top(cells_2d_23_io_fw_top),
    .io_fw_bottom(cells_2d_23_io_fw_bottom),
    .io_fw_right(cells_2d_23_io_fw_right),
    .io_sel(cells_2d_23_io_sel)
  );
  CrossBarCell cells_2d_24 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_24_io_fw_left),
    .io_fw_top(cells_2d_24_io_fw_top),
    .io_fw_bottom(cells_2d_24_io_fw_bottom),
    .io_fw_right(cells_2d_24_io_fw_right),
    .io_sel(cells_2d_24_io_sel)
  );
  CrossBarCell cells_2d_25 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_25_io_fw_left),
    .io_fw_top(cells_2d_25_io_fw_top),
    .io_fw_bottom(cells_2d_25_io_fw_bottom),
    .io_fw_right(cells_2d_25_io_fw_right),
    .io_sel(cells_2d_25_io_sel)
  );
  CrossBarCell cells_2d_26 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_26_io_fw_left),
    .io_fw_top(cells_2d_26_io_fw_top),
    .io_fw_bottom(cells_2d_26_io_fw_bottom),
    .io_fw_right(cells_2d_26_io_fw_right),
    .io_sel(cells_2d_26_io_sel)
  );
  CrossBarCell cells_2d_27 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_27_io_fw_left),
    .io_fw_top(cells_2d_27_io_fw_top),
    .io_fw_bottom(cells_2d_27_io_fw_bottom),
    .io_fw_right(cells_2d_27_io_fw_right),
    .io_sel(cells_2d_27_io_sel)
  );
  CrossBarCell cells_2d_28 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_28_io_fw_left),
    .io_fw_top(cells_2d_28_io_fw_top),
    .io_fw_bottom(cells_2d_28_io_fw_bottom),
    .io_fw_right(cells_2d_28_io_fw_right),
    .io_sel(cells_2d_28_io_sel)
  );
  CrossBarCell cells_2d_29 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_29_io_fw_left),
    .io_fw_top(cells_2d_29_io_fw_top),
    .io_fw_bottom(cells_2d_29_io_fw_bottom),
    .io_fw_right(cells_2d_29_io_fw_right),
    .io_sel(cells_2d_29_io_sel)
  );
  CrossBarCell cells_2d_30 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_30_io_fw_left),
    .io_fw_top(cells_2d_30_io_fw_top),
    .io_fw_bottom(cells_2d_30_io_fw_bottom),
    .io_fw_right(cells_2d_30_io_fw_right),
    .io_sel(cells_2d_30_io_sel)
  );
  CrossBarCell cells_2d_31 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_31_io_fw_left),
    .io_fw_top(cells_2d_31_io_fw_top),
    .io_fw_bottom(cells_2d_31_io_fw_bottom),
    .io_fw_right(cells_2d_31_io_fw_right),
    .io_sel(cells_2d_31_io_sel)
  );
  CrossBarCell cells_2d_32 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_32_io_fw_left),
    .io_fw_top(cells_2d_32_io_fw_top),
    .io_fw_bottom(cells_2d_32_io_fw_bottom),
    .io_fw_right(cells_2d_32_io_fw_right),
    .io_sel(cells_2d_32_io_sel)
  );
  CrossBarCell cells_2d_33 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_33_io_fw_left),
    .io_fw_top(cells_2d_33_io_fw_top),
    .io_fw_bottom(cells_2d_33_io_fw_bottom),
    .io_fw_right(cells_2d_33_io_fw_right),
    .io_sel(cells_2d_33_io_sel)
  );
  CrossBarCell cells_2d_34 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_34_io_fw_left),
    .io_fw_top(cells_2d_34_io_fw_top),
    .io_fw_bottom(cells_2d_34_io_fw_bottom),
    .io_fw_right(cells_2d_34_io_fw_right),
    .io_sel(cells_2d_34_io_sel)
  );
  CrossBarCell cells_2d_35 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_35_io_fw_left),
    .io_fw_top(cells_2d_35_io_fw_top),
    .io_fw_bottom(cells_2d_35_io_fw_bottom),
    .io_fw_right(cells_2d_35_io_fw_right),
    .io_sel(cells_2d_35_io_sel)
  );
  CrossBarCell cells_2d_36 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_36_io_fw_left),
    .io_fw_top(cells_2d_36_io_fw_top),
    .io_fw_bottom(cells_2d_36_io_fw_bottom),
    .io_fw_right(cells_2d_36_io_fw_right),
    .io_sel(cells_2d_36_io_sel)
  );
  CrossBarCell cells_2d_37 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_37_io_fw_left),
    .io_fw_top(cells_2d_37_io_fw_top),
    .io_fw_bottom(cells_2d_37_io_fw_bottom),
    .io_fw_right(cells_2d_37_io_fw_right),
    .io_sel(cells_2d_37_io_sel)
  );
  CrossBarCell cells_2d_38 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_38_io_fw_left),
    .io_fw_top(cells_2d_38_io_fw_top),
    .io_fw_bottom(cells_2d_38_io_fw_bottom),
    .io_fw_right(cells_2d_38_io_fw_right),
    .io_sel(cells_2d_38_io_sel)
  );
  CrossBarCell cells_2d_39 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_39_io_fw_left),
    .io_fw_top(cells_2d_39_io_fw_top),
    .io_fw_bottom(cells_2d_39_io_fw_bottom),
    .io_fw_right(cells_2d_39_io_fw_right),
    .io_sel(cells_2d_39_io_sel)
  );
  CrossBarCell cells_2d_40 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_40_io_fw_left),
    .io_fw_top(cells_2d_40_io_fw_top),
    .io_fw_bottom(cells_2d_40_io_fw_bottom),
    .io_fw_right(cells_2d_40_io_fw_right),
    .io_sel(cells_2d_40_io_sel)
  );
  CrossBarCell cells_2d_41 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_41_io_fw_left),
    .io_fw_top(cells_2d_41_io_fw_top),
    .io_fw_bottom(cells_2d_41_io_fw_bottom),
    .io_fw_right(cells_2d_41_io_fw_right),
    .io_sel(cells_2d_41_io_sel)
  );
  CrossBarCell cells_2d_42 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_42_io_fw_left),
    .io_fw_top(cells_2d_42_io_fw_top),
    .io_fw_bottom(cells_2d_42_io_fw_bottom),
    .io_fw_right(cells_2d_42_io_fw_right),
    .io_sel(cells_2d_42_io_sel)
  );
  CrossBarCell cells_2d_43 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_43_io_fw_left),
    .io_fw_top(cells_2d_43_io_fw_top),
    .io_fw_bottom(cells_2d_43_io_fw_bottom),
    .io_fw_right(cells_2d_43_io_fw_right),
    .io_sel(cells_2d_43_io_sel)
  );
  CrossBarCell cells_2d_44 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_44_io_fw_left),
    .io_fw_top(cells_2d_44_io_fw_top),
    .io_fw_bottom(cells_2d_44_io_fw_bottom),
    .io_fw_right(cells_2d_44_io_fw_right),
    .io_sel(cells_2d_44_io_sel)
  );
  CrossBarCell cells_2d_45 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_45_io_fw_left),
    .io_fw_top(cells_2d_45_io_fw_top),
    .io_fw_bottom(cells_2d_45_io_fw_bottom),
    .io_fw_right(cells_2d_45_io_fw_right),
    .io_sel(cells_2d_45_io_sel)
  );
  CrossBarCell cells_2d_46 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_46_io_fw_left),
    .io_fw_top(cells_2d_46_io_fw_top),
    .io_fw_bottom(cells_2d_46_io_fw_bottom),
    .io_fw_right(cells_2d_46_io_fw_right),
    .io_sel(cells_2d_46_io_sel)
  );
  CrossBarCell cells_2d_47 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_47_io_fw_left),
    .io_fw_top(cells_2d_47_io_fw_top),
    .io_fw_bottom(cells_2d_47_io_fw_bottom),
    .io_fw_right(cells_2d_47_io_fw_right),
    .io_sel(cells_2d_47_io_sel)
  );
  CrossBarCell cells_2d_48 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_48_io_fw_left),
    .io_fw_top(cells_2d_48_io_fw_top),
    .io_fw_bottom(cells_2d_48_io_fw_bottom),
    .io_fw_right(cells_2d_48_io_fw_right),
    .io_sel(cells_2d_48_io_sel)
  );
  CrossBarCell cells_2d_49 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_49_io_fw_left),
    .io_fw_top(cells_2d_49_io_fw_top),
    .io_fw_bottom(cells_2d_49_io_fw_bottom),
    .io_fw_right(cells_2d_49_io_fw_right),
    .io_sel(cells_2d_49_io_sel)
  );
  CrossBarCell cells_2d_50 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_50_io_fw_left),
    .io_fw_top(cells_2d_50_io_fw_top),
    .io_fw_bottom(cells_2d_50_io_fw_bottom),
    .io_fw_right(cells_2d_50_io_fw_right),
    .io_sel(cells_2d_50_io_sel)
  );
  CrossBarCell cells_2d_51 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_51_io_fw_left),
    .io_fw_top(cells_2d_51_io_fw_top),
    .io_fw_bottom(cells_2d_51_io_fw_bottom),
    .io_fw_right(cells_2d_51_io_fw_right),
    .io_sel(cells_2d_51_io_sel)
  );
  CrossBarCell cells_2d_52 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_52_io_fw_left),
    .io_fw_top(cells_2d_52_io_fw_top),
    .io_fw_bottom(cells_2d_52_io_fw_bottom),
    .io_fw_right(cells_2d_52_io_fw_right),
    .io_sel(cells_2d_52_io_sel)
  );
  CrossBarCell cells_2d_53 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_53_io_fw_left),
    .io_fw_top(cells_2d_53_io_fw_top),
    .io_fw_bottom(cells_2d_53_io_fw_bottom),
    .io_fw_right(cells_2d_53_io_fw_right),
    .io_sel(cells_2d_53_io_sel)
  );
  CrossBarCell cells_2d_54 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_54_io_fw_left),
    .io_fw_top(cells_2d_54_io_fw_top),
    .io_fw_bottom(cells_2d_54_io_fw_bottom),
    .io_fw_right(cells_2d_54_io_fw_right),
    .io_sel(cells_2d_54_io_sel)
  );
  CrossBarCell cells_2d_55 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_55_io_fw_left),
    .io_fw_top(cells_2d_55_io_fw_top),
    .io_fw_bottom(cells_2d_55_io_fw_bottom),
    .io_fw_right(cells_2d_55_io_fw_right),
    .io_sel(cells_2d_55_io_sel)
  );
  CrossBarCell cells_2d_56 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_56_io_fw_left),
    .io_fw_top(cells_2d_56_io_fw_top),
    .io_fw_bottom(cells_2d_56_io_fw_bottom),
    .io_fw_right(cells_2d_56_io_fw_right),
    .io_sel(cells_2d_56_io_sel)
  );
  CrossBarCell cells_2d_57 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_57_io_fw_left),
    .io_fw_top(cells_2d_57_io_fw_top),
    .io_fw_bottom(cells_2d_57_io_fw_bottom),
    .io_fw_right(cells_2d_57_io_fw_right),
    .io_sel(cells_2d_57_io_sel)
  );
  CrossBarCell cells_2d_58 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_58_io_fw_left),
    .io_fw_top(cells_2d_58_io_fw_top),
    .io_fw_bottom(cells_2d_58_io_fw_bottom),
    .io_fw_right(cells_2d_58_io_fw_right),
    .io_sel(cells_2d_58_io_sel)
  );
  CrossBarCell cells_2d_59 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_59_io_fw_left),
    .io_fw_top(cells_2d_59_io_fw_top),
    .io_fw_bottom(cells_2d_59_io_fw_bottom),
    .io_fw_right(cells_2d_59_io_fw_right),
    .io_sel(cells_2d_59_io_sel)
  );
  CrossBarCell cells_2d_60 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_60_io_fw_left),
    .io_fw_top(cells_2d_60_io_fw_top),
    .io_fw_bottom(cells_2d_60_io_fw_bottom),
    .io_fw_right(cells_2d_60_io_fw_right),
    .io_sel(cells_2d_60_io_sel)
  );
  CrossBarCell cells_2d_61 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_61_io_fw_left),
    .io_fw_top(cells_2d_61_io_fw_top),
    .io_fw_bottom(cells_2d_61_io_fw_bottom),
    .io_fw_right(cells_2d_61_io_fw_right),
    .io_sel(cells_2d_61_io_sel)
  );
  CrossBarCell cells_2d_62 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_62_io_fw_left),
    .io_fw_top(cells_2d_62_io_fw_top),
    .io_fw_bottom(cells_2d_62_io_fw_bottom),
    .io_fw_right(cells_2d_62_io_fw_right),
    .io_sel(cells_2d_62_io_sel)
  );
  CrossBarCell cells_2d_63 ( // @[CrossBarSwitch.scala 37:53]
    .io_fw_left(cells_2d_63_io_fw_left),
    .io_fw_top(cells_2d_63_io_fw_top),
    .io_fw_bottom(cells_2d_63_io_fw_bottom),
    .io_fw_right(cells_2d_63_io_fw_right),
    .io_sel(cells_2d_63_io_sel)
  );
  assign io_fw_bottom_0 = cells_2d_56_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_1 = cells_2d_57_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_2 = cells_2d_58_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_3 = cells_2d_59_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_4 = cells_2d_60_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_5 = cells_2d_61_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_6 = cells_2d_62_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign io_fw_bottom_7 = cells_2d_63_io_fw_bottom; // @[CrossBarSwitch.scala 77:21]
  assign cells_2d_0_io_fw_left = fw_left_reg_0; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_0_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_0_io_sel = select_onehot_0[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_1_io_fw_left = cells_2d_0_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_1_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_1_io_sel = select_onehot_1[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_2_io_fw_left = cells_2d_1_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_2_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_2_io_sel = select_onehot_2[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_3_io_fw_left = cells_2d_2_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_3_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_3_io_sel = select_onehot_3[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_4_io_fw_left = cells_2d_3_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_4_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_4_io_sel = select_onehot_4[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_5_io_fw_left = cells_2d_4_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_5_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_5_io_sel = select_onehot_5[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_6_io_fw_left = cells_2d_5_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_6_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_6_io_sel = select_onehot_6[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_7_io_fw_left = cells_2d_6_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_7_io_fw_top = 64'h0; // @[CrossBarSwitch.scala 55:28]
  assign cells_2d_7_io_sel = select_onehot_7[0]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_8_io_fw_left = fw_left_reg_1; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_8_io_fw_top = cells_2d_0_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_8_io_sel = select_onehot_0[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_9_io_fw_left = cells_2d_8_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_9_io_fw_top = cells_2d_1_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_9_io_sel = select_onehot_1[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_10_io_fw_left = cells_2d_9_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_10_io_fw_top = cells_2d_2_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_10_io_sel = select_onehot_2[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_11_io_fw_left = cells_2d_10_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_11_io_fw_top = cells_2d_3_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_11_io_sel = select_onehot_3[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_12_io_fw_left = cells_2d_11_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_12_io_fw_top = cells_2d_4_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_12_io_sel = select_onehot_4[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_13_io_fw_left = cells_2d_12_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_13_io_fw_top = cells_2d_5_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_13_io_sel = select_onehot_5[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_14_io_fw_left = cells_2d_13_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_14_io_fw_top = cells_2d_6_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_14_io_sel = select_onehot_6[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_15_io_fw_left = cells_2d_14_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_15_io_fw_top = cells_2d_7_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_15_io_sel = select_onehot_7[1]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_16_io_fw_left = fw_left_reg_2; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_16_io_fw_top = cells_2d_8_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_16_io_sel = select_onehot_0[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_17_io_fw_left = cells_2d_16_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_17_io_fw_top = cells_2d_9_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_17_io_sel = select_onehot_1[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_18_io_fw_left = cells_2d_17_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_18_io_fw_top = cells_2d_10_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_18_io_sel = select_onehot_2[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_19_io_fw_left = cells_2d_18_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_19_io_fw_top = cells_2d_11_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_19_io_sel = select_onehot_3[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_20_io_fw_left = cells_2d_19_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_20_io_fw_top = cells_2d_12_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_20_io_sel = select_onehot_4[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_21_io_fw_left = cells_2d_20_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_21_io_fw_top = cells_2d_13_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_21_io_sel = select_onehot_5[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_22_io_fw_left = cells_2d_21_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_22_io_fw_top = cells_2d_14_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_22_io_sel = select_onehot_6[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_23_io_fw_left = cells_2d_22_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_23_io_fw_top = cells_2d_15_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_23_io_sel = select_onehot_7[2]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_24_io_fw_left = fw_left_reg_3; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_24_io_fw_top = cells_2d_16_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_24_io_sel = select_onehot_0[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_25_io_fw_left = cells_2d_24_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_25_io_fw_top = cells_2d_17_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_25_io_sel = select_onehot_1[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_26_io_fw_left = cells_2d_25_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_26_io_fw_top = cells_2d_18_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_26_io_sel = select_onehot_2[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_27_io_fw_left = cells_2d_26_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_27_io_fw_top = cells_2d_19_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_27_io_sel = select_onehot_3[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_28_io_fw_left = cells_2d_27_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_28_io_fw_top = cells_2d_20_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_28_io_sel = select_onehot_4[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_29_io_fw_left = cells_2d_28_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_29_io_fw_top = cells_2d_21_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_29_io_sel = select_onehot_5[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_30_io_fw_left = cells_2d_29_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_30_io_fw_top = cells_2d_22_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_30_io_sel = select_onehot_6[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_31_io_fw_left = cells_2d_30_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_31_io_fw_top = cells_2d_23_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_31_io_sel = select_onehot_7[3]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_32_io_fw_left = fw_left_reg_4; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_32_io_fw_top = cells_2d_24_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_32_io_sel = select_onehot_0[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_33_io_fw_left = cells_2d_32_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_33_io_fw_top = cells_2d_25_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_33_io_sel = select_onehot_1[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_34_io_fw_left = cells_2d_33_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_34_io_fw_top = cells_2d_26_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_34_io_sel = select_onehot_2[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_35_io_fw_left = cells_2d_34_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_35_io_fw_top = cells_2d_27_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_35_io_sel = select_onehot_3[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_36_io_fw_left = cells_2d_35_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_36_io_fw_top = cells_2d_28_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_36_io_sel = select_onehot_4[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_37_io_fw_left = cells_2d_36_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_37_io_fw_top = cells_2d_29_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_37_io_sel = select_onehot_5[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_38_io_fw_left = cells_2d_37_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_38_io_fw_top = cells_2d_30_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_38_io_sel = select_onehot_6[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_39_io_fw_left = cells_2d_38_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_39_io_fw_top = cells_2d_31_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_39_io_sel = select_onehot_7[4]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_40_io_fw_left = fw_left_reg_5; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_40_io_fw_top = cells_2d_32_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_40_io_sel = select_onehot_0[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_41_io_fw_left = cells_2d_40_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_41_io_fw_top = cells_2d_33_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_41_io_sel = select_onehot_1[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_42_io_fw_left = cells_2d_41_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_42_io_fw_top = cells_2d_34_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_42_io_sel = select_onehot_2[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_43_io_fw_left = cells_2d_42_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_43_io_fw_top = cells_2d_35_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_43_io_sel = select_onehot_3[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_44_io_fw_left = cells_2d_43_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_44_io_fw_top = cells_2d_36_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_44_io_sel = select_onehot_4[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_45_io_fw_left = cells_2d_44_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_45_io_fw_top = cells_2d_37_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_45_io_sel = select_onehot_5[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_46_io_fw_left = cells_2d_45_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_46_io_fw_top = cells_2d_38_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_46_io_sel = select_onehot_6[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_47_io_fw_left = cells_2d_46_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_47_io_fw_top = cells_2d_39_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_47_io_sel = select_onehot_7[5]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_48_io_fw_left = fw_left_reg_6; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_48_io_fw_top = cells_2d_40_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_48_io_sel = select_onehot_0[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_49_io_fw_left = cells_2d_48_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_49_io_fw_top = cells_2d_41_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_49_io_sel = select_onehot_1[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_50_io_fw_left = cells_2d_49_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_50_io_fw_top = cells_2d_42_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_50_io_sel = select_onehot_2[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_51_io_fw_left = cells_2d_50_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_51_io_fw_top = cells_2d_43_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_51_io_sel = select_onehot_3[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_52_io_fw_left = cells_2d_51_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_52_io_fw_top = cells_2d_44_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_52_io_sel = select_onehot_4[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_53_io_fw_left = cells_2d_52_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_53_io_fw_top = cells_2d_45_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_53_io_sel = select_onehot_5[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_54_io_fw_left = cells_2d_53_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_54_io_fw_top = cells_2d_46_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_54_io_sel = select_onehot_6[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_55_io_fw_left = cells_2d_54_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_55_io_fw_top = cells_2d_47_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_55_io_sel = select_onehot_7[6]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_56_io_fw_left = fw_left_reg_7; // @[CrossBarSwitch.scala 62:29]
  assign cells_2d_56_io_fw_top = cells_2d_48_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_56_io_sel = select_onehot_0[7]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_57_io_fw_left = cells_2d_56_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_57_io_fw_top = cells_2d_49_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_57_io_sel = select_onehot_1[7]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_58_io_fw_left = cells_2d_57_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_58_io_fw_top = cells_2d_50_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_58_io_sel = select_onehot_2[7]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_59_io_fw_left = cells_2d_58_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_59_io_fw_top = cells_2d_51_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_59_io_sel = select_onehot_3[7]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_60_io_fw_left = cells_2d_59_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_60_io_fw_top = cells_2d_52_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_60_io_sel = select_onehot_4[7]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_61_io_fw_left = cells_2d_60_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_61_io_fw_top = cells_2d_53_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_61_io_sel = select_onehot_5[7]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_62_io_fw_left = cells_2d_61_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_62_io_fw_top = cells_2d_54_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_62_io_sel = select_onehot_6[7]; // @[CrossBarSwitch.scala 70:44]
  assign cells_2d_63_io_fw_left = cells_2d_62_io_fw_right; // @[CrossBarSwitch.scala 66:29]
  assign cells_2d_63_io_fw_top = cells_2d_55_io_fw_bottom; // @[CrossBarSwitch.scala 58:28]
  assign cells_2d_63_io_sel = select_onehot_7[7]; // @[CrossBarSwitch.scala 70:44]
  always @(posedge clock) begin
    fw_left_reg_0 <= io_fw_left_0; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_1 <= io_fw_left_1; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_2 <= io_fw_left_2; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_3 <= io_fw_left_3; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_4 <= io_fw_left_4; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_5 <= io_fw_left_5; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_6 <= io_fw_left_6; // @[CrossBarSwitch.scala 33:28]
    fw_left_reg_7 <= io_fw_left_7; // @[CrossBarSwitch.scala 33:28]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  fw_left_reg_0 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  fw_left_reg_1 = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  fw_left_reg_2 = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  fw_left_reg_3 = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  fw_left_reg_4 = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  fw_left_reg_5 = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  fw_left_reg_6 = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  fw_left_reg_7 = _RAND_7[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
